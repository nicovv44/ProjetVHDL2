----------------------------------------------------------------------------------
-- Company: ECE Paris
-- Engineer: Boudier Antoine - Law Nicolas - SEI group 6
-- 
-- Create Date:    17:19:00 12/25/2015 
-- Design Name: 
-- Module Name:    turret - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: Module which includes all turret components
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_STD.all;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

ENTITY turret IS
    PORT (
		clk : IN STD_LOGIC;
		reset : IN STD_LOGIC;
		posXIn_turret : IN STD_LOGIC_VECTOR (9 downto 0);
		posYIn_turret : IN STD_LOGIC_VECTOR (9 downto 0);
		beamX : IN STD_LOGIC_VECTOR (9 downto 0);
		beamY : IN STD_LOGIC_VECTOR (9 downto 0);
		beamValid : IN STD_LOGIC;
		shoot : IN STD_LOGIC;
		rotation_left : IN STD_LOGIC;
		rotation_right : IN STD_LOGIC;
		redOut_turret : OUT STD_LOGIC;
		greenOut_turret : OUT STD_LOGIC;
		blueOut_turret : OUT STD_LOGIC;
		hit : IN STD_LOGIC;
		hit_ennemy : IN STD_LOGIC;
		posXMissile : OUT STD_LOGIC_VECTOR(9 downto 0);
		posYMissile : OUT STD_LOGIC_VECTOR(9 downto 0));
END turret;

ARCHITECTURE Behavioral OF turret IS

COMPONENT missile IS
	PORT (
		clk, reset, actif, init_missile, rotation_event : IN STD_LOGIC;
		rotation: IN STD_LOGIC_VECTOR(1 downto 0);
		posXIn_missile : IN STD_LOGIC_VECTOR(9 downto 0);
		posYIn_missile : IN STD_LOGIC_VECTOR(9 downto 0);
		posXOut_missile : OUT STD_LOGIC_VECTOR(9 downto 0);
		posYOut_missile : OUT STD_LOGIC_VECTOR(9 downto 0);
		beamX : IN STD_LOGIC_VECTOR (9 downto 0);
		beamY : IN STD_LOGIC_VECTOR (9 downto 0);
		beamValid : IN STD_LOGIC;
		redOut_missile : OUT STD_LOGIC;
		greenOut_missile : OUT STD_LOGIC;
		blueOut_missile : OUT STD_LOGIC);
	END COMPONENT;	
	
TYPE image is ARRAY (natural range <>,natural range <>) OF std_logic_vector(0 to 2);
CONSTANT turret : image :=(
("111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111"),
("111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","101","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","000","111","111","111","111","110","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111"),
("111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111"),
("111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","000","111","111","111","111","111","111","110","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","100","111","111","111","111","111","111","111","111","111","111","111","000","111","111","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","111","101","111"),
("111","101","111","111","101","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","101","101","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","000","111","111","111","111","110","111","111","110","111","111","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111"),
("111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","110","110","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000"),
("111","101","111","111","111","111","111","111","111","111","111","111","111","000","111","111","100","111","111","111","110","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","110","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","100","111","111","111","111","111","111","111","111","111","111","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","000","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","101","111","111","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","100","111","111","111","111","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000"),
("111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","111","111","111","110","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","110","111","111","111","111","111","111","111","000","000","111","000","111","111","111","111","111","110","111","111","111","111","111","111","111","111","111","111","111","111","111","111","110","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","000","100","000","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000"),
("000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","000","111","111","111","111","111","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","110","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111"),
("111","000","111","111","100","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","100","111","111","111","111","111","111","111","110","111","111","111","100","000","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","111","111","111","111","111","000","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","000","000","111","000","111","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","110","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111"),
("111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","100","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","111","000","111","000","000","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","000","000","000","000","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","101","111","111","111","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111"),
("111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","111","000","111","111","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","100","111","111","111","111","111","111","111","000","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","100","000","000","000","000","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","000","000","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111"),
("111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","100","000","000","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","000","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111"),
("111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","000","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","100","100","000","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","000","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","101"),
("111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","000","111","001","111","111","111","111","111","111","111","111","111","101","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","101","111","111","101","111","111","111","111","111","111","000","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","100","100","100","100","100","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","100","111","111","100","100","100","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111"),
("111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","100","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","100","111","111","111","111","111","111","111","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","100","100","100","111","110","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","100","100","100","100","100","111","111","100","100","100","000","000","000","000","000","000","000","000","000","000","000","101","111","111","111","111","111","111","101","111","111","111","111","111","111","111","111","111","111","111","111","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","100","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111"),
("000","000","000","111","110","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","100","111","111","111","111","100","111","111","111","101","111","000","111","111","111","110","110","111","111","111","111","111","111","111","111","110","111","110","110","110","110","111","111","110","000","000","111","111","111","111","111","111","111","110","110","111","111","111","111","111","111","111","111","111","111","111","110","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","111","110","111","000","000","000","000","000","000","000","000","000","000","000","100","100","100","111","111","100","100","000","000","100","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","000","111","100","100","100","100","111","111","111","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000"),
("000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","111","111","111","100","100","000","000","111","000","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","100","100","100","100","000","000","000","000","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000"),
("000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","000","000","000","100","100","100","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111"),
("111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","100","100","000","000","000","000","000","100","100","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","100","100","100","100","111","100","111","000","111","111","111","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","011","111","111","111","111","111","111","111","000","111","111","111","111","111","111","011","111","111","111","011","111","111","111","111","111","111","011","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","011","111","111","111","111","111"),
("111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","101","111","111","111","101","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","111","111","111","000","111","000","111","100","100","100","100","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","100","100","100","100","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","101","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","101","111","111","101","111","111","111","111","111","111","111","111","111"),
("111","111","111","111","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","100","100","100","100","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","100","111","111","111","111","111","111","111","111","100","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","111","111","101","111","111","111","111","111","111","111","101","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111"),
("111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","100","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","100","111","111","111","111","111","000","000","111","111","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","100","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111"),
("111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","101","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","111","111","100","100","111","111","111","111","111","000","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","000","000","111","111","111","111","100","000","100","111","111","100","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","100","111","111","111","111","111","111","111","100","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","101","111","111","111","111","111","111","000","111","111","111"),
("111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","110","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","100","111","111","100","000","000","111","111","111","111","000","100","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","000","000","000","100","000","111","111","111","111","100","000","100","100","111","100","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","101","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111"),
("111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","100","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","110","111","111","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","000","000","000","000","000","000","000","000","000","000","100","111","100","100","000","100","111","111","111","111","000","000","100","000","000","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","000","000","000","000","000","000","111","111","000","100","000","000","100","111","100","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","100","000","000","111","111","111","111","111","111","111","111","111","111","111","110","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","110","111","111","111","111","111","111","111","111","111","111","010","111","111","111","111","111","111","000","000","111","111","111","111","111","110","111","111","111","111","111","111","010","111","111","111"),
("110","110","110","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","101","111","111","111","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","110","111","110","110","111","110","000","000","110","110","111","111","110","111","111","111","111","111","111","111","111","111","111","111","110","110","110","111","111","110","111","110","111","111","000","000","111","110","111","110","111","110","110","111","111","111","111","111","111","111","111","111","111","110","111","111","111","111","000","000","000","000","000","000","000","000","000","000","100","111","000","000","000","100","000","111","111","100","000","000","000","000","000","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","000","000","100","000","000","000","000","000","000","000","000","000","111","111","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000"),
("000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","000","000","000","000","000","000","000","000","000","000","000","000","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","000","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000"),
("000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","000","000","000","000","000","000","000","000","000","111","000","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","000","111","000","000","000","000","000","000","000","000","000","111","111","100","000","000","000","000","000","000","000","000","000","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111"),
("111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","111","111","000","000","000","000","000","000","000","000","000","111","000","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","000","111","000","000","000","000","000","000","000","000","000","111","111","111","100","000","000","000","000","000","000","000","000","111","111","111","111","000","111","111","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111"),
("111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","101","111","111","111","111","111","111","111","111","111","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","111","111","111","000","000","000","000","000","000","000","000","000","111","000","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","000","111","000","000","000","000","000","000","000","000","000","111","111","100","000","000","000","000","000","000","000","000","111","111","111","111","000","111","111","111","111","110","110","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111"),
("111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","100","111","111","000","000","000","000","000","000","000","000","000","111","000","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","000","100","000","111","111","000","000","000","000","000","000","000","111","100","100","000","000","000","000","000","000","000","000","111","111","111","111","000","111","111","111","111","111","111","111","111","011","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","011","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101"),
("111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","100","100","111","000","000","000","000","000","000","000","111","111","000","100","000","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","011","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","000","000","100","111","000","100","100","000","100","000","111","100","100","000","000","000","000","000","000","000","000","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111"),
("111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","100","100","111","000","100","000","100","100","000","111","100","100","100","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","100","000","000","100","100","100","100","000","100","100","100","000","000","000","000","000","000","000","000","111","111","111","111","000","111","011","111","111","111","111","111","111","011","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","011","111","111","111","111","111","111","111","101","111","111","111","111"),
("111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","100","100","100","100","100","100","100","100","000","000","100","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","111","111","111","100","111","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","111","111","111","111","000","111","111","111","111","111","111","111","111","011","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111"),
("111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","110","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","100","100","100","100","100","100","100","100","100","111","100","111","111","111","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","111","111","111","111","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","111","111","111","100","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001"),
("111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","111","111","111","000","000","111","111","111","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","111","111","111","111","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","111","100","100","100","111","111","111","100","100","100","100","100","000","000","100","100","100","000","000","000","000","000","000","000","111","111","110","100","000","111","111","111","111","111","111","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","111","100","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","101","111","111","000"),
("111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","111","111","111","111","010","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","100","100","100","100","100","100","100","100","100","100","111","111","110","100","100","100","111","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","111","100","100","100","100","100","100","100","100","100","100","100","000","000","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000"),
("000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","000","000","000","100","100","100","100","100","100","100","100","100","100","111","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","100","100","100","100","100","100","100","100","100","100","100","000","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","000","100","100","100","100","100","100","100","100"),
("000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","000","000","100","100","100","000","000","000","000","000","000","000","100","100","100","100","000","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","000","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","000","000","100","100","100","100","100","100","100","100","100","100","110","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","100","111","100","100","111","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","111","100","111","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","100","111","100","111","000","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100"),
("000","111","100","111","100","111","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","100","110","100","100","111","100","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","110","111","100","110","110","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","100","111","100","110","100","111","100","110","100","110","100","100","100","100","100","100","100","100","100","100","100","100","100","111","100","110","100","100","100","100","100","100","100","100","100","100","100","100","100","111","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","100","000","100","000","000","000","000","000","000","000","000","000","000","111","111","100","110","100","111","100","111","100","111","100","110","100","100","100","100","100","100","100","100","100"),
("000","111","111","100","110","100","110","100","111","100","110","100","110","100","100","100","100","100","100","100","100","100","100","100","100","100","110","100","110","100","100","100","100","100","100","100","100","100","100","100","100","100","111","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","100","000","100","000","100","100","100","000","100","000","000","000","000","000","000","000","000","000","100","000","100","100","000","000","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","100","110","110","100","111","110","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","100","111","100","100","110","111","110","100","100","100","100","100","100","100","100","111","100","000","000","000","000","000","000","111","100","111","110","111","100","111","100","110","100","110","100","111","100","111","100","111","100","100","100","100","100","111","100","111","100","110","100","111","100","111","100","111","100","100","100","100","100","111","100","111","100","110","100","111","100","110","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","100","000","000","000","000","000","111","111","110","100","110","110","110","100","111","100","111","100","110","100","111","100","111","100","111","100","100"),
("100","111","111","110","100","110","110","111","100","111","100","111","100","111","100","110","100","111","100","111","100","100","100","100","100","110","100","111","100","111","100","111","100","111","100","111","100","100","100","100","100","111","100","110","100","111","100","111","100","111","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","100","100","100","100","100","100","100","000","100","000","100","000","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","111","100","100","100","100","100","100","100","100","110","111","111","100","100","111","100","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","100","111","111","100","100","110","111","111","100","100","100","100","100","100","100","111","111","000","000","000","000","000","000","100","111","100","100","100","110","111","110","100","110","100","110","100","110","100","111","100","110","100","111","100","110","111","111","100","110","100","111","100","110","100","111","100","110","100","111","100","110","111","111","100","110","100","110","100","110","100","111","100","110","100","110","100","110","100","100","100","100","100","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","100","100","110","100","100","100","110","111","110","100","110","100","110","100","111","100","111","100","110","100"),
("000","111","100","100","110","100","100","100","110","111","111","100","110","100","110","100","110","100","110","100","111","100","111","100","111","111","111","100","110","100","111","100","111","100","110","100","111","100","111","100","110","111","111","100","110","100","110","100","111","100","110","100","111","100","110","100","100","100","100","100","100","100","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","000","100","000","000","000","000","000","000","000","000","100","111","111","100","100","100","100","100","100","100","111","111","111","100","100","110","111","100","111","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","100","100","111","100","100","100","100","100","100","100","100","100","100","100","100","111","111","111","000","000","000","000","000","111","100","111","100","111","100","110","111","110","100","111","100","110","100","110","000","111","100","110","100","110","100","111","111","110","100","111","100","111","100","111","100","111","100","110","100","110","100","110","111","110","100","111","100","110","100","110","100","110","100","111","100","111","100","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","111","110","111","000","110","100","110","100","110","111","110","100","111","100","111","100","111","100","111","100","110"),
("100","111","111","111","100","110","100","110","100","110","111","111","100","111","100","110","100","110","100","111","100","111","100","110","000","111","110","111","100","110","100","110","100","111","100","110","100","111","100","110","100","111","110","111","100","110","100","111","100","110","100","110","100","111","100","111","100","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","100","000","000","000","000","000","000","100","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","111","100","100","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","111","100","000","000","000","000","100","110","100","111","100","111","000","111","100","110","100","111","100","111","100","111","100","111","110","111","100","110","000","111","100","111","100","111","100","111","100","110","100","111","111","111","100","110","000","111","100","111","100","111","100","111","100","111","100","111","111","111","110","110","111","100","111","100","111","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","110","100","111","100","110","100","111","100","111","100","111","100","111","100","111","100","111","100","111","111"),
("000","111","111","000","111","100","111","100","111","100","111","100","111","100","111","100","111","100","110","100","111","111","111","100","111","100","111","000","111","100","111","100","111","100","111","100","111","111","111","100","111","100","111","100","111","100","111","100","111","100","110","100","111","111","111","100","111","111","100","111","100","111","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","000","100","000","000","000","000","000","000","000","100","111","111","100","100","100","100","100","100","100","100","100","100","100","100","111","100","100","100","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","011","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","111","100","100","100","100","110","100","100","100","100","100","100","100","100","100","100","100","100","111","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","100","100","100","100","100","100","100","100","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111"),
("100","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","100","100","100","100","100","100","100","100","111","111","111","111","111","111","111","111","111","111","100","100","100","000","100","100","100","000","000","000","000","000","000","000","111","100","100","100","100","100","100","100","100","100","100","100","100","110","100","100","100","100","111","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","111","000","000","000","000","000","100","100","100","100","100","000","000","000","000","000","000","000","100","000","000","000","000","100","000","100","100","000","000","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","000","000","100","100","000","100","100","100","100","000","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","000","000","000","000","000","000","000","000","000","000","100","100","100","100","100","000"),
("000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","000","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","111","100","111","100","111","000","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100"),
("100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","111","000","111","100","111","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","001","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","100","100","100","100","100","100","100","111","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","110","100","110","100","111","100","111","100","111","100","110","100","100","100","100","100","100","100","100","100","100","100","100","100","111","100","100","100","100","100","100","100","000","000","000","000","000","000","100","100","100","000","000","000","000","000","000","100","100","100","100","100","100","100","100","100","111","100","100","100","100","100","100","100","100","100","100","100"),
("100","100","100","100","100","100","100","100","100","100","111","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","111","111","000","111","100","111","100","111","100","111","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","111","100","111","100","100","100","100","000","100","000","000","000","100","000","100","000","000","000","100","000","000","000","000","000","000","000","100","000","000","000","100","000","100","000","100","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","111","100","100","100","100","100","111","100","110","100","111","100","111","100","111","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","111","111","110","100","111","111","111","100","111","100","111","100","110","100","111","100","111","100","111","100","100","100","100","100","111","100","111","100","111","100","111","100","100","100","100","000","100","100","100","100","100","100","100","000","100","000","000","000","111","100","111","100","100","100","100","100","111","100","110","100","111","100","111","100","111","100","110","100","100"),
("100","111","100","111","100","100","100","100","100","111","100","111","100","111","100","111","100","110","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","111","110","110","100","110","110","111","100","111","100","111","100","110","100","111","100","110","100","111","100","100","100","100","100","111","100","111","100","111","100","111","100","100","100","100","000","100","100","100","100","100","100","100","000","100","000","100","100","111","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","100","111","100","111","100","110","111","111","100","110","100","110","100","110","100","111","100","111","100","111","100","110","100","100","100","100","100","100","111","100","110","000","100","110","100","100","100","111","111","111","100","110","100","110","100","110","100","110","100","110","100","110","100","110","110","111","100","110","100","111","100","111","100","100","100","100","100","100","100","100","100","100","100","100","000","100","000","100","100","111","100","110","100","110","100","110","111","111","100","110","100","110","100","111","100","111","100","111","100"),
("000","100","111","100","110","100","110","100","110","111","111","100","110","100","110","100","111","100","110","100","111","100","110","100","111","100","100","100","100","111","100","111","100","111","100","100","110","100","100","100","110","111","111","100","110","100","110","100","111","100","110","100","111","100","111","100","111","110","111","100","110","100","110","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","011","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","111","100","110","100","110","100","111","110","110","100","110","100","110","100","111","100","111","100","110","100","111","100","100","111","100","100","100","100","100","100","111","110","110","100","110","100","110","100","111","111","110","100","110","100","110","100","110","100","110","100","110","100","110","100","110","111","110","100","110","100","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","100","100","111","000","111","100","110","100","110","100","110","110","110","100","111","100","111","100","111","000","111","100","110"),
("000","111","100","110","100","110","100","110","100","111","110","110","100","110","100","110","100","110","100","110","100","111","100","111","100","100","111","100","100","100","100","100","100","111","111","111","100","110","100","111","100","110","110","111","000","110","100","110","100","110","100","110","100","111","100","110","100","111","110","111","100","110","100","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","011","011","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","100","110","110","110","100","110","000","110","100","110","100","110","100","110","000","110","000","110","110","110","110","110","110","100","110","100","110","100","111","100","110","110","000","110","100","110","100","110","000","110","100","110","100","110","000","110","100","110","100","110","110","110","110","110","010","110","100","110","100","110","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","100","110","110","110","100","110","000","111","100","110","100","111","100","111","100","110","100","110","110"),
("100","111","111","100","110","110","110","100","110","100","110","100","110","100","110","100","110","100","110","100","110","110","110","100","110","111","100","110","100","110","100","111","000","111","111","100","110","100","110","100","110","100","110","000","110","000","110","100","110","100","110","100","110","111","110","100","110","100","110","100","110","110","110","100","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","000","000","000","000","011","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","111","110","110","110","110","111","110","110","110","110","110","110","110","111","110","110","110","110","110","110","110","111","110","111","111","111","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","111","110","110","110","110","110","110","110","110","110","110","111","111","111","111","110","111","111","111","110","110","110","110","110","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","111","111","110","111","110","110","110","110","110"),
("100","100","111","111","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","111","110","111","110","111","111","110","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","111","100","110","110","110","111","110","110","110","110","100","110","110","111","110","111","110","110","110","111","100","100","100","100","100","100","100","100","111","110","111","111","111","110","110","110","110","111","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","000","111","111","011","111","011","011","000","111","011","111","011","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","100","100","000","000","111","110","110","110","110","111","110","110","110","110","110","110","111","110","110","100","100","100","110","111","111","111","111","110","111","100","100","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","111","100","100","100","110","111","110","110","111","110","111","100","100","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","111","110","111","111","111","100","100","100","110","110","110","110","110","110","110","100","100","110","100","100","100","110","110","110","110"),
("100","111","100","100","100","111","111","110","110","110","110","110","110","110","110","110","110","110","110","110","111","100","100","100","110","110","110","110","110","110","110","100","100","110","100","100","100","110","111","110","110","110","110","110","110","110","110","110","110","110","110","110","111","100","100","100","110","110","110","110","110","110","110","100","100","110","111","110","110","110","110","110","110","110","110","111","110","110","110","110","110","110","111","100","100","110","110","110","110","110","110","110","111","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","000","111","111","111","000","001","111","000","011","111","011","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","100","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","110","110","110","110","110","110","110","110","110","110","110","110","110","110","111","100","100","100","110","111","110","111","110","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","111","110","110","111","100","100","100","111","110","110","110","110","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","111","110","110","111","100","100","100","110","110","110","110","110","100","100","100","100","100","100","100","100","100","110","110","110"),
("100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","111","110","110","110","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","111","111","110","110","110","100","100","100","100","100","100","100","110","110","110","110","110","110","110","000","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","111","111","111","111","111","001","001","001","011","011","011","111","011","011","011","011","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","100","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","111","100","110","100","100","100","111","111","111","111","111","100","100","100","100","100","100","100","100","100","111","110","110","110","110","110","110","110","110","110","111","110","111","100","110","100","100","100","110","111","111","110","110","100","100","100","100","100","100","100","100","100","111","110","110","110","110","110","110","110","110","110","110","110","110","100","110","100","100","100","111","111","111","111","111","100","100","100","100","100","100","100","100","100","111","110","110"),
("100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","111","110","110","100","110","100","100","100","110","110","111","110","110","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","111","110","110","100","110","100","100","100","110","110","110","110","110","100","100","100","100","100","100","100","111","110","110","110","110","110","110","110","110","110","110","110","110","100","110","100","100","100","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","000","111","111","000","000","000","000","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","110","100","111","100","100","100","100","110","100","100","110","100","100","100","100","100","100","100","100","100","110","111","110","110","110","110","110","110","110","111","111","100","110","100","111","100","100","100","100","110","100","100","110","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","110","100","111","100","100","100","100","110","100","100","110","100","100","100","100","100","100","100","100","100","110","110","110"),
("100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","110","100","110","100","100","100","100","110","100","100","111","100","100","100","100","100","100","100","100","100","111","110","110","110","110","110","110","110","111","110","110","100","110","100","110","100","100","100","100","110","100","100","111","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","111","110","100","111","100","110","100","100","100","100","110","100","100","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","000","011","111","111","111","111","111","111","011","111","111","011","111","111","011","000","011","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","100","100","100","100","100","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","100","100","100","100","100","100","100","110","110","110","110","111","110","111","100","111","110","100","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","100","111","110","100","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","110","110","111","110","110","110","100","111","110","100","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110"),
("100","100","100","100","100","100","100","110","111","111","110","110","110","110","100","110","110","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","111","111","110","110","110","110","100","110","110","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","100","110","111","100","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","100","100","100","100","100","100","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","000","001","001","111","111","111","111","111","111","011","111","011","111","111","001","000","111","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","100","100","100","111","100","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","110","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100"),
("100","100","100","100","100","100","100","100","100","110","111","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","111","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","100","100","111","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","011","111","001","111","111","111","111","111","001","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","100","100","100","100","100","100","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","100","100","100","100","100","100","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","111","111","100","100","100","100","101","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","100","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100"),
("100","100","100","100","100","100","100","100","100","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","000","000","111","111","111","111","111","000","111","111","111","111","111","111","111","111","000","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","100","100","100","100","100","100","100","100","111","111","100","100","100","100","100","100","100","000","000","000","100","100","100","100","100","100","100","000","100","100","100","100","100","100","000","000","000","000","101","101","101","100","100","100","100","101","101","101","101","101","101","101","101","101","101","101","101","101","101","101","101","101","100","100","100","100","100","000","000","000","101","100","101","100","100","101","100","100","100","100","101","101","101","101","101","101","101","101","101","100","101","101","100","100","100","100","000","000","000","000","100","100","100","100","100","100","100","100","100","100","101","100","101","101","101","101","101","101","101","101","101","101","101","101","001","101","100","100","100","100"),
("001","101","001","101","101","000","000","101","001","001","001","001","001","001","001","101","100","000","100","101","101","000","001","001","001","001","001","101","101","101","101","001","101","101","001","101","000","101","101","101","001","001","001","001","001","001","001","101","000","000","101","101","101","001","101","101","101","001","001","101","001","001","101","001","101","001","101","001","000","101","001","001","001","001","101","001","001","101","001","100","101","001","101","001","101","101","101","101","001","001","001","001","101","101","101","101","001","000","001","000","100","100","100","000","000","100","100","100","100","100","100","000","000","000","100","100","100","100","100","100","100","111","111","100","100","100","100","100","100","100","100","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","011","000","000","000","111","111","111","111","111","000","111","111","111","111","111","111","000","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","100","100","100","100","100","100","100","100","111","111","100","100","100","100","100","100","000","000","000","000","000","100","100","100","100","100","100","000","000","100","100","100","000","000","000","000","000","000","001","000","101","101","111","000","111","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","101","000","000","101","000","000","001","000","001","001","000","101","100","111","000","111","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","101","101","000","000","001","000","000","000","000","000","000","000","101","000","111","000","111","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","000","101","000","000","101","000"),
("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","111","001","111","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","111","001","111","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","111","001","011","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","100","100","100","000","000","100","100","100","100","100","000","000","000","000","000","100","100","100","100","100","100","111","111","100","100","100","100","100","100","100","100","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","000","011","000","000","000","111","111","001","111","000","000","111","111","111","111","000","000","000","111","111","011","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","100","100","100","100","100","100","100","100","100","111","100","100","100","100","100","000","000","000","000","000","000","100","100","100","100","100","100","000","100","100","100","100","000","000","000","101","000","111","000","000","001","000","111","000","110","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","011","000","011","000","001","001","000","000","010","010","000","110","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","001","000","001","000","111","001","000","000","010","111","000","111","000","000","000","001","001","001","001","001","001","001","001","001","001","000","001","000","000","000","000","000","001"),
("001","000","011","000","000","000","000","000","000","001","001","001","001","001","000","000","010","111","000","111","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","001","000","011","001","000","000","010","111","000","111","000","000","000","001","000","001","001","001","001","001","001","000","001","000","001","000","000","000","001","000","001","000","011","001","000","000","010","111","000","111","000","000","000","001","001","001","001","001","001","001","001","001","001","000","011","011","000","000","100","100","100","100","000","100","100","100","100","100","100","000","000","000","000","000","100","100","100","100","100","111","100","100","100","100","100","100","100","100","100","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","011","000","000","111","111","111","111","111","111","000","001","111","111","111","111","000","000","011","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","100","100","100","100","100","100","110","100","100","111","111","111","100","100","000","000","000","000","000","100","000","100","100","100","100","100","100","100","100","100","100","100","000","000","000","111","000","000","111","000","000","000","000","010","000","000","000","000","010","000","000","001","000","001","001","011","111","001","000","000","010","000","000","000","011","000","111","001","000","001","001","000","000","010","010","010","000","000","000","000","111","000","001","111","001","001","000","000","011","000","000","000","000","010","000","000","000","000","000","011","001","111","000","000","000","000","000","000","010","000","000","110","000","011","001","011","111","001","001","111","000","111","000","000","010","000","010","000","000","111"),
("000","000","111","010","010","000","010","000","110","010","000","000","000","010","000","000","110","010","000","010","000","000","000","000","011","011","011","001","011","011","001","000","000","000","111","000","010","000","010","010","000","000","111","000","111","010","000","000","010","000","000","010","010","000","000","010","000","000","011","000","011","111","011","000","011","011","000","000","000","000","110","000","010","000","110","110","000","000","110","010","010","000","000","000","000","011","000","001","011","000","001","001","000","001","001","000","111","011","000","000","100","100","100","100","100","100","100","100","100","100","000","100","000","000","000","000","100","100","100","111","111","111","100","100","110","100","100","100","100","100","100","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","011","011","000","000","111","111","001","111","111","111","000","111","111","111","011","111","000","000","111","011","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","100","100","100","100","100","111","111","100","100","000","000","000","100","100","100","100","100","100","100","100","100","000","000","000","000","100","100","100","100","100","100","100","000","010","000","111","000","000","111","000","000","000","000","111","000","010","010","000","010","000","000","000","000","010","000","000","111","000","000","000","000","000","000","000","000","000","111","000","000","000","001","000","000","000","000","010","000","000","010","000","110","010","000","111","000","000","000","000","111","000","000","010","000","000","000","000","010","000","000","000","000","111","000","000","000","000","000","000","000","000","010","010","000","000","000","010","111","000","000","111","000","110","000","000","110","000","010","000","000","111"),
("010","000","010","110","000","000","110","000","110","000","000","011","000","000","000","000","111","000","000","000","000","000","111","000","111","111","000","000","111","000","000","000","010","000","110","000","010","000","110","110","010","000","111","000","111","000","000","010","000","000","000","000","111","000","000","010","000","000","010","000","111","111","000","000","111","000","000","000","010","000","110","000","000","000","000","111","000","000","111","000","010","000","000","010","000","000","000","000","010","000","000","000","000","000","010","000","111","010","000","100","100","100","100","100","100","000","000","000","000","000","100","100","000","100","100","100","100","100","100","000","000","000","100","100","111","111","100","100","100","100","100","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","111","111","111","111","111","000","111","111","111","111","011","000","000","000","111","111","000","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","100","100","100","100","111","111","111","000","000","000","000","000","100","100","100","100","100","100","100","100","100","000","000","000","100","100","100","100","100","100","100","100","000","010","000","111","010","010","010","000","000","000","000","110","110","000","111","000","000","000","000","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","000","010","010","000","111","000","000","000","000","111","010","000","110","000","000","000","000","000","000","000","000","000","011","000","000","000","000","000","000","000","000","000","000","000","000","010","000","110","010","000","110","000","000","000","000","111","000","000","010","000","000"),
("000","000","000","111","000","000","110","000","010","000","000","111","000","000","000","000","010","000","000","000","000","000","010","000","111","110","000","000","111","000","000","000","000","000","010","000","010","000","010","010","010","000","111","000","010","000","000","111","000","000","000","000","010","000","000","000","000","000","010","000","111","010","000","000","000","000","000","000","000","000","010","000","000","010","000","111","000","000","111","000","000","000","000","111","000","000","010","000","010","000","000","000","000","110","000","000","111","000","000","100","100","100","100","100","100","100","000","000","000","100","100","100","100","100","100","100","100","100","100","000","000","000","000","100","111","111","111","100","100","100","100","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","011","000","000","001","111","111","111","111","111","001","111","111","011","011","111","011","111","111","111","000","011","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","100","100","100","100","111","111","100","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","100","000","100","100","100","100","100","100","100","100","110","000","000","000","010","000","010","010","000","000","000","110","110","000","111","000","000","000","000","110","000","000","000","010","010","000","000","000","000","000","000","000","010","000","000","000","000","000","000","000","000","000","000","000","010","010","000","000","000","010","000","111","010","000","000","000","110","110","000","111","000","000","010","000","010","000","000","000","010","000","000","000","000","000","000","010","000","000","000","000","010","010","010","000","010","010","000","110","000","000","000","000","111","110","000","110","000","000"),
("000","010","000","111","010","000","111","000","000","000","000","111","000","000","010","000","000","000","000","000","000","001","000","000","111","000","000","000","010","000","000","000","000","000","010","000","000","010","000","010","010","000","111","000","000","000","000","111","000","000","000","000","000","000","000","000","000","000","000","000","111","000","000","000","011","000","010","000","000","000","000","010","010","010","000","010","000","000","010","000","000","000","000","111","111","000","111","000","010","000","000","010","000","000","000","000","010","000","000","100","100","100","100","100","100","100","100","000","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","100","111","111","100","100","100","100","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","011","000","000","011","000","000","000","000","000","000","011","000","011","000","000","000","111","001","000","000","000","111","111","111","111","111","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","100","100","100","100","100","100","100","000","000","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","000","000","000","000","000","010","010","000","000","000","110","110","000","111","000","000","111","000","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","000","000","000","000","000","000","010","000","000","000","010","010","000","010","000","000","010","000","111","000","000","000","000","000","000","000","000","000","000","010","010","000","000","000","000","010","000","000","000","010","000","010","010","000","000","000","110","111","000","110","000","000"),
("000","010","000","000","111","000","010","000","000","000","000","111","110","000","110","000","000","000","000","000","000","000","000","000","110","000","000","000","000","000","000","000","000","000","000","010","000","010","000","010","110","000","110","000","000","000","000","110","111","000","111","000","000","000","000","000","000","010","000","000","111","000","000","000","000","000","010","000","000","000","000","010","010","000","000","000","010","000","010","010","000","000","000","110","111","000","111","000","000","000","000","010","000","000","010","000","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","100","100","100","100","100","100","100","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","011","000","111","011","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","000","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","010","000","010","000","111","000","000","110","000","001","000","000","111","000","111","000","000","000","000","000","000","000","111","000","000","010","000","000","000","000","000","000","110","000","010","000","010","000","000","000","111","000","000","000","000","010","000","010","000","010","000","000","111","000","010","000","000","010","000","110","000","000","000","000","000","000","000","110","000","000","000","000","000","000","000","000","111","000","000","000","000","000","000","010","000","000","000","010","111","000","111","000","000"),
("010","000","000","000","111","000","010","010","000","000","000","110","110","000","110","000","010","000","000","110","000","000","000","110","000","000","000","000","000","000","011","000","000","000","000","000","111","000","000","000","010","000","010","110","000","000","000","110","111","000","110","000","000","000","000","110","000","000","010","000","000","000","000","000","000","000","000","000","000","000","000","000","110","000","000","000","000","000","000","110","000","000","000","110","110","000","111","000","000","010","000","111","000","000","000","000","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","000","000","011","111","000","000","000","000","000","000","000","000","000","111","000","000","000","000","000","000","000","000","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","111","000","000","000","010","111","000","110","000","000","000","010","000","000","000","111","000","000","000","110","000","000","111","110","000","111","000","000","010","010","000","000","110","110","000","000","000","000","010","000","000","000","000","000","000","010","000","000","000","010","111","000","000","000","000","000","110","010","000","010","110","000","000","000","110","000","000","110","111","000","000","000","010","000","000","000","010","000","000","000","000","110","000","010","000","010","000","000","110","000","111","000","000"),
("010","000","000","000","000","000","000","010","000","000","000","010","110","000","110","000","000","010","000","110","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","000","000","000","000","000","000","010","000","000","000","000","110","000","110","000","000","010","000","111","000","110","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","000","000","000","000","111","000","010","010","010","010","000","010","000","010","000","000","010","000","111","000","000","000","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","100","100","110","100","100","100","100","100","100","100","100","100","100","100","100","100","111","111","111","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","011","000","001","011","011","000","000","000","000","000","111","111","111","011","011","111","001","011","000","000","000","000","000","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","100","100","110","111","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","000","000","000","000","000","010","111","000","000","000","000","110","000","000","000","000","111","000","000","000","111","000","000","111","110","000","000","010","110","000","110","000","000","110","110","000","000","110","111","000","010","000","000","000","111","000","000","000","000","010","010","110","000","000","000","010","010","000","000","000","000","111","000","000","000","010","000","000","110","010","000","000","110","111","000","000","010","000","000","010","000","000","000","000","000","000","111","010","000","000","010","110","000","111","000","000","000","110"),
("110","000","000","000","000","110","000","000","000","010","000","000","010","000","110","000","000","111","000","110","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","000","000","000","000","011","000","000","000","110","000","000","111","000","000","000","000","110","000","010","010","000","000","000","000","000","000","010","000","000","000","000","000","000","000","000","000","000","000","000","000","111","000","000","000","010","111","000","010","000","000","000","110","010","000","010","111","000","000","010","110","000","000","111","100","100","000","000","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","111","111","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","000","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","100","100","100","110","111","111","110","111","111","111","111","111","111","100","100","100","100","100","100","100","000","000","000","000","000","100","111","000","111","000","000","010","000","111","000","000","000","000","111","000","000","010","000","111","000","000","000","111","000","111","111","000","000","000","000","110","010","010","000","111","110","010","000","000","000","010","010","000","111","000","000","111","000","000","000","000","010","000","111","000","000","000","000","110","000","000","000","000","111","000","000","000","010","000","110","110","000","000","000","000","010","110","000","010","000","000","000","111","000","000","000","000","000","010","111","000","000","000","110","110","000","000","000","000","111"),
("000","000","000","000","000","111","000","000","000","010","111","000","010","000","000","000","010","110","000","010","110","000","000","010","111","000","000","111","111","000","000","000","000","000","000","000","000","000","000","000","000","111","000","000","000","010","111","000","010","000","000","000","110","110","000","000","111","000","000","010","110","000","000","111","010","000","000","010","000","000","000","111","000","000","000","000","000","011","111","000","000","000","110","010","000","000","000","000","111","000","000","000","111","000","000","111","110","000","000","110","100","000","000","000","000","100","100","100","100","100","100","100","100","111","111","111","111","111","111","111","111","111","111","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","011","011","000","000","000","000","000","000","000","000","111","111","111","001","000","000","000","000","000","000","000","000","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","100","100","100","100","100","100","100","000","000","000","000","000","000","110","000","000","000","000","010","000","010","000","000","000","000","010","000","000","110","000","110","000","000","000","000","000","111","010","000","000","000","010","000","110","000","000","111","000","000","000","000","000","010","110","000","010","010","000","010","000","000","000","000","110","000","110","000","000","000","000","010","000","000","110","000","110","000","000","000","000","000","110","010","000","000","000","000","010","110","000","000","010","010","000","111","000","000","000","000","010","000","111","000","000","000","000","110","000","000","111","000","111"),
("000","000","000","000","000","111","111","000","000","000","110","010","000","000","000","000","111","000","000","000","111","000","000","110","110","000","000","110","110","000","000","000","000","000","000","111","000","000","000","000","000","010","110","000","000","000","110","010","000","000","000","000","111","000","000","000","011","000","000","111","010","000","000","111","111","000","000","000","000","010","000","111","000","000","000","000","010","000","111","000","000","000","000","110","000","000","010","000","110","000","000","000","110","000","111","110","000","000","000","000","100","000","000","000","000","000","100","100","100","100","100","100","100","100","000","000","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","011","000","000","011","000","000","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","100","100","100","100","100","000","000","000","000","000","000","000","110","000","000","111","000","010","000","010","000","110","010","000","000","000","000","000","000","000","000","000","000","000","011","111","000","000","000","110","010","000","010","000","010","110","000","000","000","111","000","000","010","000","000","000","000","010","000","000","000","000","111","000","000","000","110","000","000","000","000","000","000","000","010","000","000","000","000","010","010","000","000","000","111","000","000","110","000","000","010","010","000","010","000","000","011","000","111","000","010","000","000","000","000","010","000","000","111","000","111"),
("000","010","000","000","000","000","111","000","000","000","010","010","000","000","010","000","111","000","000","000","000","000","111","010","000","000","000","000","010","010","000","000","010","010","000","111","000","000","000","000","010","000","110","000","000","000","010","111","000","000","010","000","111","000","000","000","011","000","111","010","000","000","000","000","111","000","000","000","010","111","000","110","000","000","010","000","110","000","010","000","000","010","000","110","000","000","011","000","110","000","000","000","000","000","111","010","000","000","000","000","100","000","000","000","000","100","100","100","100","100","100","100","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","011","000","001","111","000","000","000","111","000","000","000","000","000","000","111","001","000","000","000","000","000","000","000","000","000","000","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","100","100","100","100","000","000","000","000","000","000","000","110","000","000","000","000","111","000","000","111","111","000","000","000","010","000","000","000","000","000","010","000","000","010","010","000","000","010","010","000","000","110","000","010","010","000","000","111","011","000","000","111","000","000","000","000","010","010","000","000","000","111","000","000","010","111","000","000","000","010","000","000","000","000","000","010","000","000","111","010","000","000","110","010","000","000","000","000","000","000","010","000","010","000","000","010","000","111","000","000","000","010","000","000","000","000","000","010","000","010"),
("000","000","010","000","110","000","010","000","000","000","000","010","000","000","011","000","111","000","000","000","000","000","111","010","000","000","000","000","000","110","000","000","010","110","000","110","000","000","000","000","010","000","010","000","000","000","000","111","000","000","111","000","111","000","000","000","000","000","111","010","000","000","000","000","010","110","000","000","000","000","000","010","000","000","000","000","110","000","010","000","010","000","000","000","000","000","000","000","000","000","000","000","000","110","110","000","000","000","011","011","000","000","000","000","000","000","100","100","100","100","000","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","011","000","000","000","000","000","000","000","000","000","000","111","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","100","100","100","100","100","100","100","000","000","000","000","000","011","000","000","000","110","000","000","111","100","000","000","000","010","111","000","110","000","000","010","000","000","010","000","000","010","010","000","000","000","010","000","010","000","000","010","111","000","000","000","000","000","000","000","000","000","010","000","000","000","010","000","010","110","110","000","000","000","110","010","000","111","000","000","011","000","000","010","000","000","010","010","010","000","000","111","000","000","000","000","000","010","010","000","000","000","111","000","000","111","111","000","000","000","010","000","000","000","000"),
("010","000","010","000","111","000","010","010","010","010","000","000","000","000","011","000","011","000","000","000","000","010","010","000","000","000","111","010","000","010","010","000","000","010","000","110","000","000","010","000","111","000","010","000","110","010","000","000","000","000","111","000","010","000","000","000","000","010","010","010","000","000","111","010","000","110","000","000","000","000","000","010","110","000","000","000","111","000","000","110","110","000","000","000","111","000","000","000","010","000","110","000","000","111","010","000","000","111","011","000","000","000","000","000","100","100","100","100","000","100","100","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","000","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","100","100","100","100","100","100","100","000","000","000","000","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","010","010","000","110","100","000","000","000","000","000","111","000","010","010","000","110","000","000","010","000","000","010","010","000","000","000","000","000","000","000","000","010","011","000","000","000","000","000","000","000","000","000","000","010","000","000","010","000","010","110","000","000","000","000","000","111","000","010","111","000","111","000","000","000","000","000","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","000","110","010","010","000","000","000","110","110","000","110","000"),
("111","000","000","000","111","000","000","111","111","000","000","000","111","000","000","000","000","000","000","010","000","111","010","000","000","111","010","000","000","111","000","000","000","000","000","111","010","000","000","000","111","000","000","110","111","000","000","000","111","000","000","000","000","000","110","000","000","010","110","000","000","111","010","000","000","010","000","000","000","000","000","000","000","000","000","000","110","000","010","111","010","000","000","000","000","111","000","111","000","000","010","000","000","010","000","000","110","111","000","000","000","000","000","000","000","000","000","100","100","100","100","100","000","000","000","000","100","100","100","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","011","000","011","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","000","000","000","000","100","000","000","000","000","000","000","000","000","000","000","000","010","000","000","000","010","000","000","111","110","000","000","000","000","000","111","000","000","111","000","010","000","000","000","000","000","010","000","000","000","000","000","000","000","000","000","010","000","000","000","000","000","000","000","000","000","110","000","000","000","010","000","000","111","010","000","000","000","000","000","111","000","000","010","000","000","000","000","000","000","000","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","110","000","000","000","000","000","111","000","000","110"),
("000","000","000","000","111","000","110","110","110","000","000","000","110","010","000","110","000","000","111","000","000","010","000","000","010","111","000","000","000","010","000","000","000","000","000","000","010","000","000","000","110","000","010","111","110","000","000","000","010","010","000","000","000","000","110","000","000","110","000","000","010","110","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","000","110","110","000","000","000","000","000","111","000","000","010","000","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","100","100","000","000","000","000","100","100","100","100","100","100","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","011","000","000","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","111","111","111","000","000","000","000","000","000","111","000","000","111","000","010","000","000","011","000","000","000","000","000","000","000","000","000","000","000","000","110","100","000","000","100","000","000","000","100","100","100","100","000","100","100","100","000","000","000","000","000","000","000","111","010","000","110","010","000","000","010","000","000","000","000","000","000","111","000","000","000","000","000","010","010","000","000","111","000","000","000","111","000","000","000","000","010","110","000","000","000","111","000","000","000","000","000","000","010","110","000","010","010","000","000","010","000","000","000","000","000","000","111","000","000","111","000","000","110","000","000","010","010","010","000","000","111","000","000","000","000","000","000","000","000","000","000","000","010","000","000","110","010","000","000","000","000","000","111","000","000","110"),
("000","000","000","010","000","000","111","010","000","000","000","000","000","111","000","110","010","000","110","000","000","000","000","000","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","000","111","110","000","000","000","000","000","111","000","010","010","000","010","000","000","010","000","000","111","000","000","000","000","000","000","000","000","000","000","010","000","000","000","010","000","000","110","010","000","000","000","000","000","111","000","000","111","000","000","000","000","000","000","010","010","000","000","000","000","000","000","000","010","010","000","111","100","100","100","000","110","000","000","000","100","100","100","100","000","000","000","110","000","111","000","000","000","001","000","000","000","101","000","111","000","000","000","000","000","000","000","001","001","000","000","000","000","000","011","000","000","011","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","101","111","000","000","000","000","011","000","111","010","000","111","000","010","000","000","111","000","000","000","000","000","000","000","000","000","000","010","000","111","000","000","000","100","000","000","100","100","100","111","000","000","000","000","000","000","000","000","010","000","000","010","000","010","000","110","000","000","000","000","000","000","000","111","000","000","110","000","000","000","000","000","010","111","000","000","111","010","000","000","111","000","000","111","000","000","110","010","000","000","111","000","000","111","000","000","000","000","111","000","110","000","000","000","000","000","000","000","010","000","000","010","000","000","000","000","000","010","111","000","000","111","010","000","000","111","000","000","000","000","000","000","000","010","010","000","010","010","000","000","010","000","000","000","000","000","000","111","000","000","010"),
("000","000","000","010","000","000","110","000","000","000","000","000","000","111","000","000","111","000","000","000","000","000","000","000","010","000","000","000","000","000","000","000","000","000","000","010","000","000","000","010","000","000","111","000","000","000","000","000","000","111","000","000","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","110","010","000","010","010","000","000","010","000","000","000","000","000","000","111","000","000","111","000","000","111","000","000","000","110","010","000","000","111","000","000","010","000","010","010","000","111","000","000","000","000","111","010","010","010","000","000","000","000","000","000","000","000","010","111","000","000","000","000","000","000","000","000","000","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","000","000","000","000","000","000","010","010","000","111","000","000","000","000","111","110","000","110","000","000","000","000","010","000","000","000","000","000","000","000","000","000","000","000","000","100","000","110","000","000","000","000","000","000","000","000","000","010","000","010","000","010","000","010","000","000","000","000","000","000","000","111","010","000","000","000","000","000","000","010","000","010","111","000","000","111","000","000","110","000","000","111","111","000","000","111","000","000","111","000","000","111","000","000","010","000","010","000","110","000","000","000","000","000","000","000","111","110","000","000","000","000","000","000","000","000","111","110","000","000","111","000","010","111","000","000","000","110","000","000","000","000","010","000","110","000","000","000","000","000","000","010","111","000","000","010","000","000","010"),
("010","000","010","010","000","000","010","000","000","000","000","000","000","110","000","000","010","000","000","110","000","000","000","010","010","000","000","111","000","000","000","000","000","000","000","111","010","000","010","010","000","000","010","000","000","000","000","000","000","111","000","000","010","000","000","010","000","000","010","110","000","000","000","111","000","000","000","010","000","000","000","000","010","000","111","000","000","000","000","000","000","000","010","000","000","011","000","000","010","000","000","110","010","000","000","010","111","000","000","111","000","000","000","000","010","010","000","111","000","000","000","000","010","010","010","011","000","000","000","010","010","000","010","000","000","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","000","000","000","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","000","000","000","111","000","000","000","010","000","000","000","010","000","010","010","000","000","000","110","111","000","110","000","000","000","000","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","000","000","000","010","000","000","000","000","000","000","000","110","111","000","000","000","000","010","000","111","000","000","111","000","000","111","000","010","110","000","000","000","111","000","000","010","000","110","010","000","000","010","000","000","010","000","000","000","110","000","000","000","000","000","000","000","111","111","000","000","000","000","111","000","111","000","000","111","000","000","111","000","110","010","000","000","010","110","000","000","010","000","010","000","111","000","000","000","000","000","000","000","111","010","000","000","000","000","010"),
("111","000","010","000","000","000","000","000","000","000","111","000","000","010","000","000","000","000","000","000","111","000","000","111","110","000","000","111","000","000","000","111","000","000","000","000","010","000","010","000","000","000","000","000","000","000","010","000","000","010","000","000","010","000","000","000","111","000","000","110","111","000","010","111","000","000","010","111","000","000","000","000","010","000","111","000","000","000","000","000","000","000","111","011","000","000","000","000","000","000","010","000","111","111","000","000","111","000","010","111","000","000","000","000","000","010","000","110","110","000","000","000","010","111","000","111","000","000","000","000","010","000","000","111","000","000","000","000","000","000","000","000","000","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","011","000","000","000","111","111","001","111","101","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","101","111","001","000","000","111","000","000","000","011","000","000","000","000","000","000","110","000","000","000","000","110","000","110","000","000","010","010","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","000","010","000","000","000","000","000","000","000","000","000","000","010","110","000","000","000","111","110","000","010","000","000","010","000","000","110","000","010","010","000","000","000","010","000","000","010","000","010","000","000","000","000","000","000","110","110","000","000","000","000","000","110","000","000","000","000","000","111","000","000","000","010","111","000","111","000","000","010","000","000","110","000","110","000","000","000","010","010","000","000","110","000","000","000","010","000","000","000","000","000","000","000","110","111","000","000","000","000","110"),
("010","000","010","000","000","000","000","000","000","000","111","000","000","000","000","000","010","000","010","000","111","111","000","000","111","000","000","111","000","000","000","111","000","000","010","000","010","000","010","000","000","000","000","000","000","000","111","111","000","000","000","000","000","000","010","000","111","110","000","000","111","000","010","110","000","000","110","010","000","000","111","000","000","000","010","000","000","000","000","000","000","000","011","111","000","000","000","000","110","000","111","000","000","010","000","000","110","000","000","010","000","111","000","000","000","000","000","000","110","000","000","000","010","111","000","110","000","000","110","000","110","000","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","000","000","000","111","111","000","111","111","111","111","001","111","001","000","000","000","000","000","000","000","000","000","000","000","000","001","111","111","111","111","111","001","000","000","000","000","000","000","011","000","000","000","000","010","000","010","000","110","000","000","110","000","010","000","000","010","000","111","000","000","000","000","000","000","000","001","000","000","010","000","000","000","000","000","000","111","000","000","000","000","000","010","000","010","000","111","000","000","000","000","000","111","010","000","000","000","000","010","000","000","000","111","000","000","000","000","000","000","000","000","010","010","000","000","000","000","000","000","000","000","010","110","000","000","000","000","000","000","000","110","111","000","000","000","000","000","111","000","000","000","000","000","010","000","000","000","111","000","000","000","000","000","000","000","010","000","010","000","000","000","000","010","000","000","000","111","010","000","000","000","000","000","000","010","000","010","000","000","111","000","000","000","111","111"),
("000","000","010","000","000","000","000","000","000","000","111","111","000","000","000","000","111","000","110","000","000","111","000","000","111","000","110","010","000","000","111","000","000","000","111","000","000","000","010","000","000","000","000","000","000","000","000","111","000","000","000","000","111","000","110","000","000","111","000","000","111","000","010","010","000","000","010","000","000","000","111","000","000","000","000","000","000","000","000","010","000","000","000","111","000","000","000","110","111","000","010","000","000","010","000","000","111","000","010","000","000","010","000","000","000","000","110","000","110","000","110","000","000","010","000","000","000","000","111","000","111","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","000","010","000","110","000","000","000","010","000","000","000","000","111","111","000","111","000","111","111","111","111","111","011","000","000","000","000","000","000","000","000","000","001","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","111","000","000","000","110","111","000","010","000","010","000","110","010","000","111","111","000","000","000","010","000","000","111","011","000","011","000","000","000","111","000","000","111","010","000","000","000","010","010","000","000","000","111","000","000","000","000","111","111","000","000","010","010","000","000","000","000","000","111","000","000","000","010","000","000","000","000","000","010","000","000","000","000","000","000","000","000","000","010","000","000","000","000","000","010","000","000","110","000","000","000","000","111","111","000","000","000","010","000","000","000","000","000","010","000","000","000","110","000","000","000","000","000","010","000","000","000","000","000","000","000","010","111","111","000","000","000","000","000","111","010","000","000","000","000","010","000","000","000","111","000"),
("000","000","000","000","000","000","000","000","000","000","000","111","000","000","000","111","010","000","110","000","000","010","000","000","010","000","010","000","000","000","010","000","000","000","111","010","000","000","000","000","000","000","000","110","000","000","010","111","000","000","000","111","010","000","111","000","000","010","000","000","111","000","010","000","000","000","000","000","000","010","110","111","000","000","000","000","000","111","110","000","000","000","000","011","000","000","000","111","000","000","000","000","000","000","000","000","000","110","000","000","000","000","000","000","000","000","111","000","000","000","010","111","000","010","000","000","000","110","010","000","111","110","000","000","000","111","000","000","111","010","000","010","000","000","000","000","000","000","111","010","000","000","000","110","010","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","111","111","111","000","000","111","000","000","000","000","000","000","000","000","000","000","000","000","000","010","111","000","000","000","111","010","000","000","000","000","111","000","000","000","111","000","000","111","110","000","000","110","111","000","010","000","000","111","110","000","000","010","111","000","010","000","000","000","111","000","000","000","010","000","000","111","010","000","010","000","000","110","010","000","000","000","000","010","000","000","000","111","000","000","111","110","000","000","000","000","000","000","000","000","110","110","000","000","000","000","000","010","010","000","000","000","000","111","000","000","111","000","000","111","000","000","010","110","000","000","000","000","010","000","000","000","110","000","000","010","110","000","000","000","000","010","000","000","000","010","000","000","000","000","000","000","000","111","010","000","000","000","110","000","000","000","000","000","111","000"),
("000","000","000","000","000","111","010","000","000","000","000","110","000","000","000","111","010","000","010","000","000","000","000","000","000","010","000","010","000","000","000","000","000","010","010","111","000","000","000","000","000","111","110","000","000","000","000","010","000","000","000","111","010","000","000","000","000","000","000","000","000","110","000","000","000","000","000","000","000","000","000","110","000","000","000","000","010","111","000","000","000","110","000","000","000","000","000","110","000","000","000","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","110","110","000","010","000","010","010","000","000","000","000","111","000","000","000","011","000","010","110","110","000","000","000","111","000","111","000","000","111","111","000","000","110","111","000","000","000","000","000","111","000","000","000","000","000","000","000","000","000","000","111","000","000","111","111","111","000","000","000","000","000","111","000","000","111","111","111","000","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","010","000","110","000","000","000","010","110","000","000","000","000","111","000","000","000","010","000","110","110","000","000","000","000","111","010","010","000","010","111","000","000","000","000","110","110","000","110","010","000","111","000","110","000","000","000","000","010","000","000","110","010","000","000","111","000","000","000","000","000","000","010","000","000","010","000","000","111","110","000","010","010","000","011","010","000","010","111","110","000","010","010","000","111","000","000","000","010","000","000","000","000","111","000","000","010","110","000","010","111","000","010","000","000","000","000","010","000","000","000","000","000","111","010","010","110","000","000","010","000","000","000","010","000","000","010","000","000","010","000","000","010","000","000","110","110","000","000","000","000","010","000"),
("010","000","000","000","111","111","000","000","000","010","000","000","000","000","000","110","010","000","000","110","000","000","000","000","000","000","000","000","000","000","000","000","010","000","000","110","000","000","000","000","111","111","000","000","000","110","000","000","000","000","000","010","000","000","000","110","000","000","000","000","000","000","000","000","000","000","000","010","000","010","000","000","110","000","000","000","111","000","000","000","000","111","110","000","000","000","000","000","000","000","000","111","000","000","010","110","000","000","000","000","000","000","010","000","000","000","000","111","000","010","000","010","010","000","000","000","000","111","000","000","000","010","000","111","110","000","000","000","000","110","000","010","000","111","010","000","000","000","000","010","000","000","111","000","000","111","000","000","000","000","000","000","000","000","000","000","000","000","000","111","000","000","000","000","111","000","000","111","111","000","000","000","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","000","010","000","000","000","000","110","000","000","111","000","111","000","000","000","000","000","111","010","000","000","000","000","010","110","000","000","111","010","000","000","000","000","010","110","000","010","110","000","110","000","000","000","000","000","000","010","000","000","000","111","000","000","010","000","010","000","010","000","000","111","000","000","010","000","000","010","111","000","000","111","000","000","000","000","000","010","111","000","000","111","000","010","000","111","000","010","000","000","000","000","111","000","000","000","110","000","000","110","000","110","000","010","000","000","111","000","000","110","000","000","010","111","000","000","110","010","000","000","010","000","000","000","000","000","000","000","111","000","000","000","000","000","000","111","000","000","000","000","000","000"),
("000","000","000","000","111","000","000","000","000","111","010","000","000","000","000","000","000","000","000","010","000","000","110","000","000","000","000","000","000","110","000","010","000","000","000","000","000","000","000","110","110","000","000","000","010","110","010","000","000","000","000","000","000","000","000","010","000","000","000","111","000","000","000","000","000","010","000","010","000","000","010","000","000","000","000","111","010","000","110","010","000","010","111","000","000","000","000","000","000","010","000","000","000","000","000","111","010","000","010","010","000","000","000","010","000","010","000","010","000","000","000","111","000","000","111","000","110","000","000","010","000","010","000","010","010","000","000","000","000","000","110","000","111","111","000","000","010","000","000","000","110","000","111","000","000","000","010","000","000","111","000","111","000","000","000","000","000","000","000","000","111","000","000","000","111","000","000","111","001","000","000","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","111","000","010","000","010","010","000","000","000","000","000","000","111","000","000","000","000","010","010","000","000","000","111","110","000","000","000","000","111","000","000","000","110","010","000","010","000","000","000","000","110","010","000","111","000","000","000","111","000","000","000","110","000","000","000","000","110","000","111","000","000","010","111","000","000","000","000","000","110","000","000","110","010","000","000","000","000","000","111","000","000","111","010","000","000","010","010","010","110","000","000","000","010","000","000","000","010","000","000","000","000","111","000","111","000","000","111","111","000","000","000","000","000","111","000","000","010","010","000","000","000","111","000","010","000","000","000","000","111","000","000","000","110","000","000","110","000","111","000","000","000","000"),
("000","000","000","111","000","000","010","000","000","000","111","000","000","000","000","000","000","110","000","000","010","000","000","110","010","000","010","000","000","010","000","110","000","000","000","000","000","000","000","110","000","000","110","000","000","010","111","000","000","000","000","000","000","010","000","000","010","000","000","111","110","000","110","000","000","111","000","000","111","000","110","000","000","000","000","111","000","000","010","010","000","000","110","000","010","000","010","000","000","111","000","000","000","000","000","010","111","000","000","110","000","000","000","000","000","111","000","010","000","010","000","111","010","000","111","000","000","000","000","111","000","000","110","000","000","000","000","000","000","010","000","000","110","000","000","000","000","000","000","000","000","000","111","000","000","000","000","000","000","000","000","111","000","000","000","000","000","000","000","000","111","111","111","000","111","111","000","111","000","111","111","111","111","000","000","000","000","000","000","000","111","000","000","111","000","010","000","000","010","000","000","010","010","000","000","000","000","000","000","000","000","111","000","000","000","010","000","000","000","000","000","111","111","000","000","000","000","000","000","000","000","000","000","000","010","000","000","000","000","010","010","000","111","000","000","000","000","000","000","010","010","000","110","010","110","110","000","111","000","000","000","111","010","000","000","000","000","010","000","000","000","010","000","000","000","000","000","110","000","000","000","010","000","000","000","000","000","111","000","000","000","000","000","000","010","110","000","010","000","010","010","000","111","000","000","000","111","010","000","000","000","000","111","000","000","000","010","000","000","000","000","111","000","010","000","000","000","011","000","000","000","010","000","000","000","000","111","000","111","000","000"),
("000","000","000","111","000","000","010","010","000","000","111","000","000","000","010","000","000","111","000","000","110","000","000","111","110","000","010","111","000","000","000","000","111","000","110","000","000","000","000","010","000","000","000","111","000","000","111","000","010","000","010","000","000","111","000","000","010","000","000","000","111","000","010","111","000","000","000","000","000","111","000","110","000","000","000","010","000","000","000","010","000","000","010","000","111","000","010","000","000","010","111","000","000","000","000","000","111","000","000","110","010","010","000","000","000","111","000","000","000","110","000","000","110","000","110","000","000","000","000","111","110","000","111","000","000","000","000","000","000","000","000","000","111","000","000","000","000","000","000","000","010","000","010","000","000","000","000","000","011","000","000","000","110","000","000","000","000","000","000","000","111","000","000","111","000","000","000","001","111","000","000","000","000","000","000","000","000","000","000","010","110","000","000","111","000","000","000","000","111","000","000","010","000","000","000","000","000","000","010","000","000","111","000","000","000","010","000","000","000","000","000","110","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","000","000","000","000","000","111","000","000","010","010","000","111","000","000","000","000","000","000","000","010","000","000","000","000","000","000","000","000","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","000","000","000","000","000","110","000","000","000","110","000","111","000","000","000","010","000","000","010","111","000","000","000","000","010","000","000","000","011","000","000","000","000","010","000","111","000","000","000","000","000","010","000","010","000","010","000","110","110","000","010","000","000"),
("000","000","000","000","000","000","000","110","000","000","010","000","110","000","110","000","000","010","111","000","000","000","000","000","110","000","000","110","010","000","000","000","000","111","000","111","000","000","000","111","000","000","000","110","000","000","010","010","111","000","010","000","000","010","111","000","000","000","000","000","111","000","000","111","010","000","010","000","000","111","000","111","000","000","000","000","000","000","000","010","000","000","000","110","111","000","010","000","000","000","111","010","000","000","000","000","111","000","000","010","010","010","000","000","000","111","000","000","000","000","000","000","010","000","010","010","000","000","000","110","110","000","111","000","000","000","000","010","000","000","010","000","000","000","000","000","000","000","000","000","010","000","000","000","000","000","000","000","000","000","000","000","000","010","000","000","000","000","000","000","000","000","000","000","000","111","000","000","000","000","000","000","000","000","000","000","000","000","111","000","110","110","000","110","000","000","000","000","110","010","000","110","000","000","000","000","000","000","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","110","000","000","010","110","000","110","000","000","000","000","000","000","000","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","110","000","000","010","110","000","111","000","000","000","111","000","000","000","110","000","000","000","000","000","000","011","000","000","000","011","000","000","000","000","010","000","000","000","000","000","010","000","010","000","110","000","111","010","000","000","000","000"),
("000","000","000","000","000","000","000","110","000","010","010","110","111","000","010","000","000","000","111","000","000","000","000","000","111","000","000","000","110","000","010","000","000","010","000","111","000","000","000","000","000","110","000","110","000","010","000","010","111","000","010","000","000","000","111","010","000","000","000","000","111","000","000","000","010","000","000","000","000","000","000","110","000","000","000","000","000","110","000","010","000","110","000","110","010","000","000","010","000","000","010","111","000","000","000","000","010","000","000","000","010","000","000","000","000","010","000","110","111","000","000","000","000","000","010","010","000","000","000","010","110","000","010","000","000","010","000","111","000","000","000","000","000","000","000","000","000","000","000","010","000","000","000","000","000","000","000","000","000","000","000","000","000","110","000","000","000","000","000","000","000","000","000","000","000","111","000","000","000","000","000","000","000","000","000","000","000","111","000","000","000","010","000","010","010","000","000","000","110","111","000","111","000","010","000","000","010","000","000","010","000","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","011","000","000","000","000","000","000","111","000","000","000","010","000","111","010","000","000","111","110","000","111","000","000","000","010","000","000","000","010","000","010","000","000","000","000","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","000","111","010","000","000","010","111","000","111","000","000","000","110","000","000","000","111","000","010","000","000","000","000","111","000","000","000","000","000","000","000","000","010","000","000","000","000","000","111","000","111","000","110","000","111","000","000","000","010","000","000","000")
);

signal destruction : std_logic := '0';
signal sennemydown : std_logic;
									
signal newPosX_turret : std_logic_vector(10 downto 0);
signal newPosY_turret : std_logic_vector(10 downto 0);
signal sigValid_turret, romSig_turret : std_logic;

signal sposXCurrent_turret : std_logic_vector(9 downto 0);
signal sposYCurrent_turret :  std_logic_vector(9 downto 0);

signal sred_turret : std_logic;
signal sblue_turret : std_logic;
signal sgreen_turret : std_logic;

signal sredOut_turret: std_logic;
signal sblueOut_turret : std_logic;
signal sgreenOut_turret : std_logic;

signal reg1_turret : std_logic_vector(31 downto 0):= x"00000000";
signal mux1_turret : std_logic_vector(31 downto 0):= x"00000000";
signal comp_turret : std_logic;

signal actif : std_logic;
signal init_missile : std_logic;

signal srotation_missile : std_logic_vector(1 downto 0);
signal rotary_event : std_logic;

signal sposXInit_missile : std_logic_vector(9 downto 0) := "0100111000";
signal sposYInit_missile : std_logic_vector(9 downto 0) := "0110010000";
signal sposXIn_missile : std_logic_vector(9 downto 0);
signal sposYIn_missile : std_logic_vector(9 downto 0);
signal sposXOut_missile : std_logic_vector(9 downto 0);
signal sposYOut_missile : std_logic_vector(9 downto 0);

signal sred_missile : std_logic;
signal sblue_missile : std_logic;
signal sgreen_missile : std_logic;

BEGIN

	destruction <= hit or destruction when rising_edge(clk);
	sennemydown <= hit_ennemy when rising_edge(clk);

	--INPUT PART

	rotary_event <= '1' when rotation_left = '1' or rotation_right = '1'
		else '0' when srotation_missile = "01" or srotation_missile = "10";

	actif <= '0' when sennemydown = '1'
		else '1' when shoot = '1' -- when button is pushed, actif = '1'
			else '0' when(sposYIn_missile = "0000000000" and shoot = '0');
			
	init_missile <= '1' when actif = '1' --  initialization of a missile 
		else '0' when sposYIn_missile = "0110001111"; -- posYMissileInit - 1

	--

	--SYNCHRONISATION PART
			
	--reg1_turret is equal to mux1 when rising edge
	reg1_turret <= (others => '0') when reset='1' 
		else mux1_turret when rising_edge(clk);

	--comp is equal '1' when reg1_turret = defined value
	comp_turret <= '1' when reg1_turret = x"0003FF81" --reg1_turret = x"02FAF081" --50M = 1s
		else '0';		

	-- timer 	
	mux1_turret <= std_logic_vector(unsigned(reg1_turret) + 1) when  comp_turret = '0'
		else (others => '0');

	--

	--MISSILE PART

	missile_function : missile port map (
		clk => clk,
		reset => reset,
		actif => actif,
		init_missile => init_missile,
		rotation_event => rotary_event,
		rotation => srotation_missile,
		posXIn_missile => sposXIn_missile,
		posYIn_missile => sposYIn_missile,
		posXOut_missile => sposXOut_missile,
		posYOut_missile => sposYOut_missile,
		beamX => beamX,
		beamY => beamY,
		beamValid => beamValid,
		redOut_missile => sred_missile,
		greenOut_missile => sgreen_missile,
		blueOut_missile => sblue_missile);

	posXMissile <= sposXOut_missile;
	posYMissile <= sposYOut_missile;	

	srotation_missile <= "01" when rotation_left = '0' and rotation_right = '1'
		else "10" when rotation_left = '1' and rotation_right = '0'
			else "00";

	sposXIn_missile <= (others => '0') when reset = '1'
		else sposXOut_missile when comp_turret = '1'
			else sposXInit_missile when init_missile = '1' or sposYIn_missile = "0000000000";

	sposYIn_missile <= (others => '0') when reset='1'
		else sposYOut_missile when comp_turret = '1'
			else sposYInit_missile when init_missile = '1' or sposYIn_missile = "0000000000";

	--

	--DISPLAY PART

	sposXCurrent_turret <= (others => '0') when reset='1'
		else posXIn_turret;

	sposYCurrent_turret <= (others => '0') when reset='1'
		else posYIn_turret;

	newPosX_turret <= std_logic_vector(('0'&unsigned(beamX))-('0'&unsigned(sposXCurrent_turret)));
	newPosY_turret <= std_logic_vector(('0'&unsigned(beamY))-('0'&unsigned(sposYCurrent_turret)));

	sigValid_turret <= '0' when destruction = '1'
						else '1' when signed(newPosX_turret)<331 and signed(newPosX_turret)>=0 and signed(newPosY_turret)>=0 and signed(newPosY_turret)<95 and beamValid='1' 
							else '0';

	sred_turret <= '1' when (turret((to_integer(unsigned(newPosY_turret(6 downto 0)))),(to_integer(unsigned(newPosX_turret(8 downto 0))))) = "100"
						or turret((to_integer(unsigned(newPosY_turret(6 downto 0)))),(to_integer(unsigned(newPosX_turret(8 downto 0))))) = "110"
						or turret((to_integer(unsigned(newPosY_turret(6 downto 0)))),(to_integer(unsigned(newPosX_turret(8 downto 0))))) = "101"
						or turret((to_integer(unsigned(newPosY_turret(6 downto 0)))),(to_integer(unsigned(newPosX_turret(8 downto 0))))) = "111")
						else '0';
						
	sgreen_turret <= '1' when (turret((to_integer(unsigned(newPosY_turret(6 downto 0)))),(to_integer(unsigned(newPosX_turret(8 downto 0))))) = "010"
						or turret((to_integer(unsigned(newPosY_turret(6 downto 0)))),(to_integer(unsigned(newPosX_turret(8 downto 0))))) = "110"
						or turret((to_integer(unsigned(newPosY_turret(6 downto 0)))),(to_integer(unsigned(newPosX_turret(8 downto 0))))) = "011"
						or turret((to_integer(unsigned(newPosY_turret(6 downto 0)))),(to_integer(unsigned(newPosX_turret(8 downto 0))))) = "111")
						else '0';
						
	sblue_turret <= '1' when (turret((to_integer(unsigned(newPosY_turret(6 downto 0)))),(to_integer(unsigned(newPosX_turret(8 downto 0))))) = "001"
						or turret((to_integer(unsigned(newPosY_turret(6 downto 0)))),(to_integer(unsigned(newPosX_turret(8 downto 0))))) = "101"
						or turret((to_integer(unsigned(newPosY_turret(6 downto 0)))),(to_integer(unsigned(newPosX_turret(8 downto 0))))) = "011"
						or turret((to_integer(unsigned(newPosY_turret(6 downto 0)))),(to_integer(unsigned(newPosX_turret(8 downto 0))))) = "111")
						else '0';
							
	romSig_turret <= '1' when ((sred_turret = '1' or sblue_turret = '1' or sgreen_turret = '1') and sigValid_turret = '1') 
		else '0';
					
	sredOut_turret <= '1' when (sred_turret = '1' and romSig_turret = '1') 
		else '0';
		
	sgreenOut_turret <= '1' when (sgreen_turret = '1' and romSig_turret = '1') 
		else '0';

	sblueOut_turret <= '1' when (sblue_turret = '1' and romSig_turret = '1')
		else '0';

	redOut_turret <= sredOut_turret or sred_missile;	
	greenOut_turret <= sgreenOut_turret or sgreen_missile;	
	blueOut_turret <= sblueOut_turret or sblue_missile;				

	--

END Behavioral;