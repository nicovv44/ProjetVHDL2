----------------------------------------------------------------------------------
-- Company: ECE Paris
-- Engineer: Boudier Antoine - Law Nicolas - SEI group 6
-- 
-- Create Date:    17:25:12 12/25/2015 
-- Design Name: 
-- Module Name:    end_game - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: Module which includes all end game components
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity end_game is
	PORT(
		isTurretHit : IN STD_LOGIC;
		ennemy1Down : IN STD_LOGIC;
		ennemy2Down : IN STD_LOGIC;
		ennemy3Down : IN STD_LOGIC;
		beamX : IN STD_LOGIC_VECTOR (9 downto 0);
		beamY : IN STD_LOGIC_VECTOR (9 downto 0);
		beamValid : IN STD_LOGIC;
		rOUT, gOUT, bOUT : OUT STD_LOGIC);
END end_game;

architecture Behavioral of end_game is

TYPE imageV is ARRAY (0 to 75) OF std_logic_vector(0 to 221);
TYPE imageL is ARRAY (0 to 92) OF std_logic_vector(0 to 399);
	
signal looseImg : imageL :=(
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000111111111111111000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000001111111111111110001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111110011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000011111111111111000111111111111100000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000001111111111111100011111111111111100000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111100111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000111111111111110001111111111111111111100000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000011111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000001111111111111000111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110001111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000111111111111100011111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110001111111111101111111100000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000001111111111111000111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000011111111111100111111000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000111111111111100111111111111111100000011111111111111100111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100111111111111111110111000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000111111111111011111111111111110000000001111111111110000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110001111111111111111110000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000011111111111001111111111111111000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100011111111111111111100000000000000000001111111111000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000111111111100111111111111111110000000000000000000000000111110000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000111111111111111110000000000000000000000111111111100000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000001111111110001111111111111110000000000000000000000000001111110000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110001111111111111111000000011100000000000000111111111110000000000000111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000011111111100011111111111111100000000000000000000000000011111100000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100001111111111111110000110011111000000000000011111111111000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000111111110000111111111111100000111111000000000000011100111111000000000000000000000000000000000000000001111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000011111111111111000011110011111111000000000001111111111100000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000001111111110001111111111111000011111111110000000111111011111111000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000111111111111000000111110011111111100000000000111111111110001111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000111111111000011111111111000000011111111111111111111101111111110000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000111111111100000001111100111111111111000000000011111111111111111111111100000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000"),
("0000001111111110000011111111100000000011111111111111111111111111111100000000000000000000000000000000000000001111111111000111111111110000000000000000000000000111110000000000000000000000000000000000000000000000000000000000111111111111000001111111111000000011111100111111111111000000000011111111111111111111111000011111111111111111000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000011111111100000111111110000000000011111111100011111101111111111000000000000000000000000000000000000000001111111100000011111111111111111111100000000000111111111100000000000000000000111111111110000000000000000000000000111111111110000011111100000000000011111100011111111111100000000001111111111111111111100011111111111111111111000000000000000000000000000000000000000000000000000000111100000000000000"),
("0000011111111000000111111100000000000011111111110111111011111111110000000000000000000000000000000000000000001111111000000001111111111111111111111111110011111111111110000000000011111111111111111111110000000000000000000001111111111100000011111000001100000011111100011100111111110000000001111111111111111111000011111111111111111110000000000000000000000000000000000000001111111000001111111111110000000000"),
("0000111111110000001111110000110000000011111111111111110111111111000000000000000000000000000000000000000000001111110000000000111111111111111111111111111111111111111111001111111111111111111111111111111000000000000000000011111111110000000111111111111100000011111100011000011111110000000000111111111111111111000111111111111111111100000000000000001111111111000000000000111111111111111111111111111000000000"),
("0001111111100000001111110011110000000011111111111111111111111110000000000000000000000000000000000000000000011111000000000000111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111111110000000111111111111100000011111100011000001111111000000000011111111111111110001111111111111111110000000000000011111111111111110000000111111111111111111111111111111000000000"),
("0001111110000000001111111111110000000011111011111111111111111100000000000000000000000000000000000000000000001111100000000000111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111100000001111111111111100000011111100111100001111111100000000001111111111111000011111111111110000000000000001111111111111111111111111111111111111111111111111111111111100000000"),
("0011111100000000001111111111110000000011111001111110111111111000000000000000000000000000000000000000000000001111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111000000001111111111111100000011111100111100001111111110000000000111111111110000111111111111000000000000011111111111111111111111111111111111111111111111111111100111111110000000"),
("0011111100000000001111111111110000000111111001111101111111111000000000000000000000000000000000000000000000001111111100000000011111111111110011111111111111111110011111111111111111111111111111000111111111000000000000000111111111000000001111111111111100000011111100111110001111111110000000000011111111100001111111111100000000000111111111111111111111110001111111111111110000001111111111000111111110000000"),
("0011111100000000001111111111110000000111111001111001111111111000000000000000000000000000000000000000000000001111111110000000011111111111000001111111111111111000001111111111111111111111111100000011111111100000000000001111111110000000001111111111111000000011111100111111111111111111000000000011111110000011111111111000000111111111111111111111111111000000111111111111100000000111111111000011111111000000"),
("0011111100000000001111111111110000000111111001110011111111111111000000000000000000000000000000000000000000000111111110000000011111111110000000111111111111100000000111111111111111111111100000000001111111110000000000001111111110000000001111111111111000000011111100111111111111111111000000000001111110000111111111100000111111111111111111111111110000000000011111111111000000000011111110000011111111100000"),
("0011111000000000001111111111110000000111111000100111111111111111000000000000000011111000000000000000111000000011111110000000011111111000000000001111111111000000000001111111111111110000001100000000111111110000000000001111111100000000001111111111111000000001111100111111111111111111000000000001111100001111111111100011111111111111111111111100000011000000001111111110000000000011111100000001111111110000"),
("0111111000000000001111111111110000000111111000011111111111111111110000000001111111111110000000000011111100000011111110000000011111100000000000000111111100000000000000000011111100000000001111000000011111111000000000011111111100000000001111100111111000000001111100000000111111111000000000000001111100001111111111111111111111111111111110000000000111110000000111111100000000000001111000000000000111110000"),
("0111111000000000001111111111110000000111111000000000000111111111111110111111111111111111100000001111111111000111111110000000011110000111100000000011111001100000000000000111111100000000011111100000001111111100000000001111111100000000001111100111111000000001111100000000000110000000000000000001111000001111111111111111111111111111111111000000000111110000000011111011000000000000111000000000000011110000"),
("0111111000000000011111100111110000000011111000111111111000111111111111111111111111111111111001111111111111111111111110000000011000011111110000000011100111111000000000001111111110000000011111110000000111111110000000001111111000000000001111000011111000000001111100111111111111111111000000000001111000001111111111111111111111111111111111100000000111111100000001111111110000000000101100000000000111111000"),
("0111111000000000011111100111110000000011100001111111111100000111111111111111111111111111111111111111111111111111111111000000000001111111110000000000000111111100000000011111111111000000011111111000000011111110000000001111111000000000001111000011111000000011111100111111111111111111000000000001110000001111111111111111111111111111111111110000001111111110000000111111110000000000011110000000001111111000"),
("0111111000000000111111000111110000000011001001111111111110000000111111111111111111111111111111111110011111111111111111000000000011111111110000000000011111111110000000011111111111000000111101111100000001111110000000001111111000000000001111000011111000000011111100011111111111111111100000000011110000001111111111111111110011111111111111110000001111111111000000011111111000000000111111111111111111111100"),
("0111111000000000111111000011110000000000110011111111111111000000001111111111111111111111111111111100001111111111111111000000001111111111110000000000011111111110000000111111111111000000111000111100000000111110000000000111111000000000001111000011111000000011111100011111111111111111100000000011110000001111111111111110000000111111111111110000001111011111000000001111111100000000111111111111111111111100"),
("0111111000000000111111000011110000000001110011111110001111100000000011111111110000001111111111110000000111111111111111000000011111111111110000000001111111111110000000111111111111000000111000111110000011111110000000000111111000000000001111000011111000000011111110011111111111111111100000000011110000001111111111110000000000001111111111110000001111011111100000111111111100000000111111111111111111111100"),
("0111111000000000111111000011110000000011111001111110001111110000000001111111110000000111111111000000000011111111111111100000011111111111110000000001111111011110000000111111111111000000111001111110000111111110000000000111111000000000011111000011111000000011111110011111110001111111100000000011110000000111111111100000000000000011111111110000001111111111100001111111111100000001111111111111111111111100"),
("0011111000000000111110000011100000000111111001111111001111111000000000111111100000000111111000000000000001111111111111100000011111110111110000000001111110011110000000111110001111000000111111111110001111111100000000000011111000000000011111000011111000000011111110011111110001111111100000000011111000000001111111010000000000000000011111110000001111111111100111111111111100000001111111111111111111111100"),
("0011111000000000111110000011100000000111111001111111111111111000000000111111110000000111110000000000000000001111111111100000011111100111111000000011111110011110000000111110001111000000111111111110111111111100000000000011111000000000011111000011111000000011111110011111110001111111100000000011111000000000111111111100000000000000111111110000001111111111101111111111111100000001111111111111111111000000"),
("0011111000000000111110000011100000000011111001111111111111111000000000011111111000000000011111000000000000111111111111100000011111100011111000000011111100011110000000111110001111100000111111111001111111111000000000000011111000000000011111000011111000000011111110011111110000111111100000000111111100000000111111111111000000000000111111111000001111111111011111111111111100000001111111111100000000000000"),
("0011111100000001111110000011100000000011111000001111111111111000000000001111111100000000111111110000000001111111111111100000011111000011111000000011111100011110000000111110000111100000111111110011111111111000000000000011111000000000011111000011111000000001111110011111111111111111100000000111111100000000111111111111100000000011111111110000001111111100111111111111111100000001111111111000000000000000"),
("0011111100000001111110000011100000000011111000000000000000000000000000001111111111111111111111111100000011111111111111100000011111000011111000000011111100001110000000111110000111000000011111001111111111110000000000000011111000000000011111000111111000000001111110001111111111111111100000000111111110000000111111111111111000000011111111110000000111100111111111100011111100000001111111110000000000000000"),
("0011111100000001111110000111100000000011111001111100000000111100000000011111111111111111111111111100000011111111111111100000011111000011111000000011111100001110000000111100000111000000010000111111111111110000000000000011111100000000011111000111111000000001111110001111111111111111100000000111111110000000011111111111111000000011111111110000000100001111111111000011111100000001111111110000000000000000"),
("0011111100000000111110000111100000000011111000111111111111111100000000011111110111111111111111111100000011111111111111100000011111000011111000000011111100001110000000111100000111000000001111111111111111100000000000000001111100000000011111000111111000000001111110001111111111111111000000000111111110000000011111111111111000000011111111110000000011111111111100000011111100000001111111100000000000000000"),
("0011111100000000111111000011100000000011111000111111111111111100000000111111000011111111111111111100000011111110111111100000011111000011111000000011111100001110000000111100000111000000011111111111111111000000000000000001111100000000011111101111111100000001111110000000110001111111000000000111111100000000011111100111111000000011111111110000000111111111111000000111111100000001111111100000000000000000"),
("0001111110000000111111000111100000000011111000111110000111111100000000111111000011111111111111110000000011111100111111100000011111000011111000000011111100001110000000111100000111000000111111111111111110000000000000000001111100000000001111111111111100000001111100001111111111000010000000000111111100000000011111000111111000000011111111110000001111111111100000000111111000000011111111100000000000000000"),
("0000111110000000111111000111100000000011111000111110000011111100000000111110000011111111111111111000000011111100111111100000011111000011111000000011111100001110000000111100000111000000111111111111111100000000000000000001111100000000001111111111111100000001111100011111111111111000000000001111111100000000011111000011111000000011111111110000001111111111000000001111111000000011111111100000000000000000"),
("0000111111000000111111000111100000000011111000111111000011111100000000111110000111110001111111111100000011111000011111000000011111000011111000000011111100001110000000111100000111000000111111111111111000000000000000000000111110000000001111111111111100000011111100011111111111111100000000001111111100000000011110000011111000000011111111110000001111111110000000001111111000000011111111100000000000000000"),
("0000011111000000111111000111100000000111111000111111111111111100000000111110001111000111111111111100000011111000011111000000011111000011111000000011111100001110000000111110000111000000111111111111110000000000000000000000111110000000001111111111111100000011111100011111111111111110000000011111111100000000011110000011111000000011111111110000001111111000000000011111111000000011111111100000000000000000"),
("0000011111100000011111111111100000000111111100111111111111111100000000011110011110001111111111111100000011111000011111000000011111000011111000000011111100011110000000111110000111000000111111111111100000000000000000000000111111000000000111111111111100000011111100111111111111111110000000011111111110000000111110000011111000000011111111110000001111110000000001111111111000000011111111100000000000000000"),
("0000001111100000011111111111100000000111111101111100001111111100000000011110011110011111111111111100000011111000011111000000011111000011111000000011111100011110000000111110000111000000111111111111000000001111100000000000111111100000000111111111111000000011111000111111111111111110000000111111111110000000111110000011111000000011111111110000001111110000000111111111111000000011111111110000000000000000"),
("0000001111110000001111111111100000001111111101100000000000111100000000011110111100111111111111111100000011111000011111000000011111000011111000000011111110011110000000111110000111000000111111111111111111111111111000000000011111110000000111111111111000000011111000111111001111111110000001111111111111000000111110000011111000000011111111110000001111110000011111111111111000000011111111110000000000000000"),
("0000000111111000001111111111100000011111111100000011111000001000000000011111111100111111100001111100000011111000011111000000011111100111111000000011111111111110000000111111000111000000111111111111111111111111111000000000011111111000000011111111111000000011111000111111000111111100000011111111111111000000111110000011111000000011111111110000001111110000111111111111111000000011111111111000000000000000"),
("0000000011111100000011111111100000111111111100111111111111100000000000011111111000111111000001111100000011111000111111000000011111110111111000000011111111111110000000111111101111000000111111111111111111111011111000000000011111111100000011111111110000000011111000111110001111111100000111111111111111000000111110000011111000000111111111110000001111111111111111111110111000000011111111111110000000000000"),
("0000000011111110000011111111100001111111111101111111111111110000000000111111111000111110000001111000000011111000111111000000011111111111111000000011111111111110000000111111111111000000111111111111111111100001110000000000001111111110000001111111110000000111111000111110011111111000001111111111111111000000111110000011111000000111111111110000001111111111111111111000011000000011111111111111000000000000"),
("0000000011111111000000111111000011111100111101111111111111100000000001111111110000111100000001111000000011111000111111000000011111111111111000000011111111111110000000111111111111000000111111111111111110000111110000000000001111111111000000011111100000001111111000111111111111110000011111111111111111000000111110000011111000000111111111110000001111111111111111110001111000000011111111111111100000000000"),
("0000000001111111100000011111001111111000111101111111111111000000000011111111110000111100000001111000000011111101111111000000011111111111111000000011111111111110000000111111111111000000111111111111111100001111100000000000000111111111100000001111000000001110111000111111111111100000111111111111111111000000111110000011111000000111111111110000001111111111111111000011111000000011111111111111111000000000"),
("0000000000111111110000000111111111111001111101111111111111000000000111111111100000111100000011111000000011111111111111000000011111111111111000000111111111111110000000111111111111000000111111111111110000111111000000000000000111111111110000000111000000111100111100111111111111000001111111111111111111000000111110000011111000000111111111110000000111111111111100001111111000000001111111111111111111000000"),
("0000000000011111111100000001111111111011111001111111111110000000011111111111100000111100000011111000000011111111111111000000011111111111111100000011111111111110000000111111111111000000001111111111100011111111000000000000000011111111111000000011110111111100111100111111111110000011111111111111111111000000111110000011111000000111111111110000000011111111111000111111111000000001111111111111111111100000"),
("0000000000001111111111000000011111111111111001111111111100000000111111111111000000111100000011111000000011111111111111000000011111111111111000000011111111111110000000111111111111000000000001111111000111111100000000000000000011111111111100000000111111111111111100111111111100000111111111111111111111000000111110000011111000000111111111110000000000011111110001111111000000000000111111111111111111100000"),
("0000000000001111111111110000001111111111111001111111110000000011111111111111000000111100000011111000000011111111111110000000011111111111110000000000110001111110000000111111111110000000000000011100011111111100000000000000000011111111111110000000011111111111111100111111111000001111111111111111111111000000111111000011111000000111111111100000000000000111000111111110000000000000011111111111111111000000"),
("0000000000000111111111111111100001111111111001111100000000001111111111111110000000111100000111111000000011111111111110000000001111111111000000000000000011111110000000111111111000000000000000000000111111110000000000000000000001111111111111100000000011111111111100111111110000111111111111111111111111000000111111000111111000000111111110000000000000000000011111111000011000000000000000111111111110000000"),
("0000000000000001111111111111111111011111110001110000001111111111111111111110000000111110011111111000000011111111111110000000000111111111100000000000001111111110000000011111111011111000000000000011111111100000000000000000000000111111111111110000000000000001111100011111100011111111111111111111111111000000111111111111111000000111111110111100000000000000111111111101111110000000000001111111111100000000"),
("0000000000000000111111111111111111111111110000000111111111111111111111111100000001111111111111110000000011111111111100000000000011111111110000000011111111111110000000011111111111111100000000000111111111000000000000000000000000011111111111111110000000000000000000000000111111111111111111111111111111000000111111111111111000000111111111111111000000000001111111111111111111000000000111111111111000000000"),
("0000000000000000011111111111111111111111111111111111111111111111111111111100000000111111111111110000000001111111110000000000000001001111111000000111111111111110000000001100111111111111000000001111111110000000000000000000000000001111111111111111111000000000000000000111111111111111111111111111111111000000111111111111111000000111111111111111110000000111111111111111111111100000001111111111110000000000"),
("0000000000000000001111111111111111111111111111111111111111111111100111111100000000111111111111110000000001111111000000000000000000111111111111111111111111111110000000001000111111111111110000111111111100000000000000000000000000000001111111111111111111111111111111111111111111111111110000111111111110000000111111111111111000000011111111111111111000001111111111111111111111110000011111111111000000000000"),
("0000000000000000000111111111111111111111111111111111111111111110000011111000000000111111111111100000000001111111011110000000000001111111111111111111111111111110000000000001111111111111111001111111110000000000000000000000000000000000000001111111111111111111111111111111111111111111100000011111111110000000011111111111111000000011111111111111111110011111111111111111111111111000111111111110000000000000"),
("0000000000000000000000001111111111111111111111111111111100000000000011111000000000001111111100000000000001111111111111100000000011111111111111111111111111111111000000000001111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111111111101100000000011111111100000000000001111111110000000001111111111111111111111111111111111111111111111111111111111000000000000000"),
("0000000000000000000000000000111011111111100010001111000000000000000011111000000000000111111000111000000000111111111111110000000111111111111111111111111111111111000000000011111111111111111111111110000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000011111111000000000000000011111000000000001111111111111111111111111111111111100111111111111111111100000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000111111100000000111111111111111000011111111111111111111111111000111111110000000111111111111111111111110000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000011111111110000000000000000000111111111111111111110001111111111111111110000000001111111111111111100000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000001111100000000000000001111111100000000011111111111111111111111111111111111111111000000000111111111100000000000000111111111000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000011111111111110000000000000111111111111111111110000000001111111111111000000000000011111111111111000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000001111110000000000000011111111110000000001111111111111111111111110011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000011111111111111111111000000000000000111111000000000000000011111111111100000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000111111000000000000111111111111000000000111111111111111111110000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000111111111111111111000000000000000000001100000000000000000000111111110000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000011111100000000011111111111111100000000000011111111111111100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000011111111111111111100000000000000000000000000000000000000000000000100000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000001111111100000111111111111111110000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111100000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000")
);


signal winImg : imageV :=(
"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"000000001111110000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"000000111111111100000000000000000000000000000001000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"000001111111111111000000000000000000000000000111100000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"000011111111111111100000000000000000000000011111110000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"000011111111111111110000000000000000000001111111110000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"000111111111111111111000000000000000000111111111111000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"000111111111111111111000000000000000011111111111111000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"001110000001111111111100000000000001111000111111111100000000000000111000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"001110000000111111111100000000000111100000011111111100000000000000110000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"001100000000011111111110000000011110000000011111111100000000000000100000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"001100000000001111111110000001111100000000011111111110000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"001000000000001111111111000111100000000000001111111110000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"001000000000000111111111011111000000000000001111111110000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"000000000000000011111111111100000000000000000111111111000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"000000000000000011111111110000000000000000000111111111000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"000000000000000011111111100000000000000000000111111111000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"000000000000000001111111100000000000000000000011111111000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"000000000000000001111111100000000000000000000011111111000000000010000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000001000000000000000000000000000001110000000000000001100000",
"000000000000000001111111100000000000000000000011111111000000000111000000000000000000000001111000000000000001111111111111111100000000000000001111000000000000000000000011100000000000110000000000000011111000000000000011110000",
"000000000000000001111111100000000000000000000011111111100000001111100000000000000000000011111110000000000011111111111111111100000000000000011111110000000000000000001111110000000011111000000000000111111100000000001111110000",
"000000000000000000111111110000000000000000000011111111100000111111111000000000000000000111111111100000000111111111111111111100000000000000111111111100000000000000011111111000000111111100000000011111111110000000011111111000",
"000000000000000000111111110000000000000000000001111111100001111111111100000000000000001111111111111000000111111111111111111100000000000011111111111111000000000000111111111100001111111110000000111111111110000000111111111000",
"000000000000000000111111110000000000000000000011111111000011111111111110000000000000111111111111111110000111111111111111111100000000001111111111111111111000000001111111111100011111111111000001111111111110000001111111111100",
"000000000000000000111111110000000000000000000011111111000011111111111110000000000001111111111111111100000000111111110000000000000000111111111111111111111110000011111111111110111111111111000011111111111111000011111111111100",
"000000000000000000111111110000000000000000001111111111000000111111111100000000000111111111111111111000000000111111110000000000000011111111001111111111111111000110011111111111100111111111100010000111111111001111111111111110",
"000000000000000000111111111111100000000011111111111111000000111111111000000000111111111110111111111000000000111111110000000000000011111111000011111111111111000000001111111111000011111111000000000111111111011100011111111110",
"000000000000000000111111111111111111111111111011111111000000111111111000000000111111111110001111110000000000111111110000000000000011111111000000111111111111000000001111111110000001111110000000000111111111111000011111111110",
"000000000000000000111111111000111111111111000011111111000000111111111000000000001111111110000011110000000000111111110000000000000011111111000000000111111111000000001111111110000000111100000000000111111111110000001111111110",
"000000000000000000111111110000000000000000000011111111000000011111111000000000000111111110000000100000000000111111110000000000000011111111000000000111111111000000001111111110000000111000000000000111111111100000001111111110",
"000000000000000000111111110000000000000000000011111111000000111111111000000000000111111110000000000000000000111111110000000000000011111111000000000111111111000000001111111110000000010000000000000111111111000000001111111111",
"000000000011111100011111110000000000000000000011111110000000111111111000000000000111111110000000000000000000111111110000000000000011111111000000000111111111000000001111111110000000000000000000000111111111000000000111111111",
"000000001111111110111111110000000000000000000011111110000000111111111000000000000111111110000000000000000000111111110000000000000011111111000000000111111111000000001111111110000000000000000000000111111111000000000111111111",
"000000011111111111111111110000000000000000000011111100000000111111111000000000000111111110000000000000000000111111110000000000000011111111000000000111111111000000001111111110000000000000000000000111111111000000000111111111",
"000000111111111111111111110000000000000000000111111100000000111111111000000000000111111110000000000000000000111111110000000000000011111111000000000111111111000000001111111110000000000000000000000111111111000000000111111111",
"000000110000111111111111110000000000000000000111111100000000111111111000000000000111111110000000000000000000111111110000000000000011111111000000000111111111000000001111111110000000000000000000000111111111000000000111111110",
"000000000000001111111111110000000000000000000111111000000000111111111000000000000111111110000000000000000000111111110000000000000011111111000000000111111111000000001111111110000000000000000000000111111111000000000111111110",
"000000000000000111111111100111111111000000001111111000000000111111111000000000000111111110000000000000000000111111110000000000000011111111000000000111111111000000001111111110000000000000000000000111111111000000000111111110",
"000000000000000011111111111111111111111100001111110000000000111111111000000000000111111110000000000000000000111111110000000000000011111111000000000111111111000000001111111110000000000000000000000111111111000000000111111110",
"000000000000000011111111111100000111111111001111110000000000111111111000000000000111111110000000000000000000111111110000000000000011111111000000000111111111000000001111111110000000000000000000000111111111000000000111111100",
"000000000000000001111111100000000000000111111111100000000000111111111000000000000111111110000000000000000000111111110000000000000011111111000000000111111111000000001111111110000000000000000000000111111111000000000111111100",
"000000000000000001111111000000000000000000111111000000000000111111111000000000000111111110000000000000000000111111110000000000000011111111000000000111111111000000001111111110000000000000000000000111111111000000001111111100",
"000000000000000001111111000000000000000000111111000000000000111111111000000000000111111110000000000000000000111111110000000000000011111111000000000111111111000000001111111110000000000000000000000111111111000000001111111000",
"000000000000000000111111000000000000000000111110000000000000111111111000000000000111111110000000000000000000111111110000000000000011111111000000000111111111000000001111111110000000000000000000000111111111000000001111110000",
"000000000000000000111110000000000000000001111110000000000000111111111000000000000111111110000000000000000000111111110000000000000011111111000000000111111111000000001111111110000000000000000000000111111111000000011111110000",
"000000000000000000111110000000000000000001111100000000000000111111111000000000000111111110000000000000000000111111110000000000000011111111000000000111111111000000001111111110000000000000000000000111111111000000011111100000",
"000000000000000001111100000000000000000011111000000000000000111111111000000000000111111110000000000000000000111111110000000000000011111111000000000111111111000000001111111110000000000000000000000111111111000000111111000000",
"000000000000000001111100000000000000000011110000000000000000111111111000000000000111111110000000000000000000111111110000000000000011111111000000000111111111000000001111111110000000000000000000000111111111000000111110000000",
"000000000000000001111000000000000000000011110000000000000000011111111000000000000111111110000000000000000000111111110000000000000011111111000000000111111111000000001111111110000000000000000000000111111111000001111100000000",
"000000000000000001111000000000000000000111100000000000000000111111111000000000000111111110000000000000000000111111110000000000000011111111000000000111111111000000001111111110000000000000000000000111111111000011111000000000",
"000000000000000011110000000000000000001111000000000000000000111111111000000000000111111110000000000000000000111111110000000000000011111111000000000111111111000000001111111110000000000000000000000111111111000111110000000000",
"000000000000000011100000000000000000001110000000000000000000111111111000000000000111111110000000000000000000111111111000000000000111111111100000000111111111000000001111111110000000000000000000000111111111001111000000000000",
"000000000000000011100000000000000000011100000000000000000000111111111000000000000111111110000000000000000001111111111000000000000111111111111000000111111111000000011111111110000000000000000000000111111111011110000000000000",
"000000000000000111000000111111111100111000000000000000000001111111111000000000001111111111100000000010000001111111111110000100001111111111111110000111111111000000011111111111000000110000000000000111111111111000000000000000",
"000000000000000111000011111111111111110000000000000000000011111111111100010000001111111111111100000110000111111111111111011100001111111111111111110111111111000000111111111111110011100000000000001111111111100000000000000000",
"000000000000001110001111111111111111100000000000000000000011111111111111110000011111111111111111001100000111111111111111111000001111111111111111111111111110000001111111111111111111000000000000001111111111000000000000000000",
"000000000000001100111111111111111111000000000000000000000000111111111111100000011111111111111111110000000000111111111111110000000000011111111111111111111000000000001111111111111110000000000000011111111100000000000000000000",
"000000000000011111111111111111111110000000000000000000000000011111111110000000001111111111111111100000000000001111111111000000000000000011111111111111000000000000000011111111111000000000000000011111110000000000000000000000",
"000000000000011111111111111111111100000000000000000000000000001111111100000000000000111111111111000000000000000011111110000000000000000000111111111100000000000000000000111111110000000000000000111111000000000000000000000000",
"000000000000111110000000000111111000000000000000000000000000000111111000000000000000000111111110000000000000000001111100000000000000000000001111111000000000000000000000011111100000000000000000111100000000000000000000000000",
"000000000000110000000000000001110000000000000000000000000000000011110000000000000000000001111000000000000000000000111000000000000000000000000111100000000000000000000000001111000000000000000000111000000000000000000000000000",
"000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000001110000000000000000000000000000",
"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000",
"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000",
"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000",
"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000",
"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000",
"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000001100000000000000",
"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000111110000000000000",
"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000001111100000000000000",
"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000111111100000000000000",
"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000",
"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000",
"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
);

signal win, loose : std_logic;
signal newPosX : std_logic_vector(10 downto 0);
signal newPosY : std_logic_vector(10 downto 0);
signal sigvalid : std_logic;
signal romsig : std_logic;
signal posXCurrent : std_logic_vector(9 downto 0);
signal posYCurrent : std_logic_vector(9 downto 0);

BEGIN

	posYCurrent <= "0011010111";
	posXCurrent <= "0001111000" when loose = '1'
							else "0011010000" when win = '1'
								else "0000000000";
	win <= (not isTurretHit) and ennemy1Down and ennemy2Down and ennemy3Down;

	loose <= isTurretHit;

	newPosX <= std_logic_vector(signed(std_logic_vector(('0'&unsigned(beamX))))-(signed(posXCurrent)));
	newPosY <= std_logic_vector(signed(std_logic_vector(('0'&unsigned(beamY))))-(signed(posYCurrent)));
	sigValid <= '1' when signed(newPosX)<222 and signed(newPosX)>=0 and signed(newPosY)>=0 and signed(newPosY)<76 and beamValid='1' and win='1'
		else '1' when signed(newPosX)<400 and signed(newPosX)>=0 and signed(newPosY)>=0 and signed(newPosY)<93 and beamValid='1' and loose='1'
		else '0';
	romSig <= '1' when (winImg(to_integer(unsigned(newPosY(6 downto 0))))(to_integer(unsigned(newPosX(8 downto 0))))='1' and sigValid='1' and win='1')
		else '1' when (looseImg(to_integer(unsigned(newPosY(6 downto 0))))(to_integer(unsigned(newPosX(8 downto 0))))='1' and sigValid='1' and loose='1')
		else '0';

	rOut <= 	'1' when (loose='1' and romSig='1')
					else '0';

	gOut <= 	'1' when (win='1' and romSig='1') 
					else '0';

	bOut <= 	'0';
	
END Behavioral;